// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:51:51 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Wu6vFupNggAK7oOaFUjX346Uar7rygtQIUD2O7VdfCEapn6ROnfhoPPmG9q9DayE
s7NpnJOp4TXr2uQGLmxoGhxzY8tvWgr6Mr0Q3KgS19Ied1E7gvEJ1pIcLdHZl6Lr
bH86CiOnSoqkcXUiJasgGTYB4d5M+lgQfULx0GdlW9E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11040)
z+23Cpn73+GXQGIzQlwoxnp1oofj6ADYpfjb4YZENCk92dEdppivDkAKLf57kxp9
51iKwT7uT0oof2nLd/8Z8dUmJavi/SPck84u93swHCoUpW4volvJnZFFGeoa2zdU
NTn5kbgFJFbMvMTtbuMZ/lp/23jLZRcmVELbneXu0sc3mcdycFu7blTrApzl5YP7
c3XGjjJgFM0QvyJFz9cH9MQ58eB3ydiqiLSvoAW/zy8++CSZt7Pm4iGs2VJpq3mM
QAmAOEC0PUZq9yHk1mnvXYTYYvMa7iEC7UsG0MiiFuvMIRU4rYoWEbw4TOAEobPT
IHyrLLKFKluwoY/7NkAJMzmL24+jnJA55xhz3i4qmDi8tjSeJGwedlEOW3cUvJ77
u5gcJJRSajV1Vngpy9w1vCQreS9j5zAR29Jw4e5TLEacFWqTJNQ5hDvCRa71MA5k
SjdLMt64W+/D9JH28Jdj3vN6JgFCbmfNMUm63vjhVVy7OeOJZpShJ/i1Z5i/4XfE
4t9c86na2V8dHhSLIaQLv1lZoROU4thwXnwei2EKW2odwFHeTsy/fQUBWcFCq7z1
VTnkRejcwtvEF/NRVDzpRRJd+D4OQCV6/dTOQSGVhDaxg01NTx5NY5zS2/l97N8a
zpzKMaA0stvcu9uFfwQN4Cf5aR2OESB5qWMEUAr6VADWp8E3Vd8oRliyJxHFPFDh
QsshmGLTOsbmfvFxlPJlb+YqPcrhpdC6uSyqloomKGT3Ik8fb9vR2Vp0a/PkBbes
4ecfI6fhXP/P9vHb4YbgPzh8zicN7MqyDxGLHaenSJ4vfFJIjOLcfTMP8+FbuAsd
YkwN5IS37tTiHRDfDCCUMU+IdFxcljFnHTJ8ELYm4k6fMhYwzZMx+Ry0Dwdql5lz
/tYpszeMkjAMCl0f0kEG8CXKC0qNUL83HZCMSLj0ZRYGkC2pisDPcTb6Ie7ghhhJ
zmC36kfJ1f7mJ3v7fs093TpRcdak/eyOhr2sYTVmJh7rpAlNfON8t3LI7IoXvsAI
JJ5ru+shFTgPSD2INKyFByTMPeRZKayVUvum8XahkmTm1ML3rVDeJ39MlbKawYSV
vh58uf/TSfM1mByQtH453fyRRyzoquDYrhjbZaM1jy4X7qvKIR6hol+eqZ2j2kAR
Xnjywb9mA0JM5q8cN7zPkS4i1lof1AFmkeD/97ESbmIATwCSv2TNuBU0mQozNW0H
DTFVJ1xU0XQLXX4DPsysfRRSNHOxx9wedDht784MUo8dvX4VyGoh4CDfTMaVadac
dMwFi+OXbc3XT1evRC6O4Z19LvFE/aPjyyEfbTmBD+syZHQKhyLNjPyaldK+Jo2K
46TKWfZEQLbbJgc/gR5i4esyMlvMrcklTW2U0i3nBMTEvb/3PTYoJzdz3m1O+YOg
kAZiXQrsjlVQCZSIVYT7EkNbzr8W8t5qN1Iv7RjK5WQiiV6HVw9/qR07KZU/lLgs
O5rbj/+0/EOiJ7wkklXYx1fyaMqT3ltoHWDuJ5Dp/TGlXI7E2oeo4y7kH6pRreq6
D1NOrFoiQaAeijn5roNo04+t0Fcpjbm95V/HwGIpFSWJQH03nTjniZ0CGWDUNRzX
tN2GAjHVXpBDzUwszqJamlGpYstVXR5U4YpiR0zHjLbFZ9QsmhHkaClJMLBoyfMj
/uh9Yhn892aU/fL3jkMR0HihPCi+mv+/icgXcdmU31ASNQsvQwD6nvsRx/UkQt4k
T8Mm9ByqJUJ1+mTgAcGobIGabSzpJpLsRgcqslJrm7sXJ1Y7WPqeTBz5WTjAUaJx
M40neI5+kgTKq4JPps3vimuNyOsecZ75g4iY2jLEApdaj1Ps6pdxsXB3trwbxUpi
sluvJuD4yHOA52zSb16ECtkoVFJ3B7j8cweuEjMSxUYn9Yz9DL/Q3kmQdOvYOkGt
LdHWfHGc1QAdABAdgwK6d2sULx18G8j8fHbEU07SfZ+E8Al4pN0uVarKXYX7QcNz
4FqIa5sKhe+yUcFUGV39oc8nXyYmDvffYzOmgyA8kpqb8XSB0CY7JXyf0LA/imQ/
Vtp+O1Ox94IJwHvP9bh5cVPhhlwms+mShzfwdzdgoNZBpSt0P1ZxXQ3udc013Xcy
yjuMqBB/OzkVhDoFZuHZ6Cc5D6teEt7ozvDprZRCmvoxEvlb0LZ1a2Fy6aHoq7pa
OKrFrxJEEii1HTrDPOk7Urg/JKijfNVZU8FWogN/iP4AdS+WmgMNUOFyL9LGGQBP
MKtRhiy5YSTK8wTrVqlSfOpf2g7Wni5E/aroq0C9QWdaPRDFPjaQwiJ4hadKuCOE
GBjkgRhtDmDGwNaZJuWc2HIlOkjJ8T6X1joZHh5U2EJ88Fh7nyGlGcplfAQwvGbI
Euc+Oub3JySdzeFyymr9PvlNOW5dMCMlJ64V1o1tRT4kn03bWZS96MXWqRd3NmTN
txR1PZhZ6po6OsXZDpxw7Da1DbTCo5Q+dmT7F/T6tEGn885mJaLPnLL5JhX2mEHq
eBC3w87/m4wT3FLjiYmaUaZO/M9xIqoXU+Rk3BRAWnwr49hpmtRbjCnD30BTOsf7
U9RLtv5gnzGwgsiifN3WKl00aV+8Alrfw1g565+n7ncp+R6ZRsTPSdVnD1IbPFWC
eMuPFjktmbYmT7oW+PsrbYgQVN/ny6tARBdinM5zDz56oy16Ew5y/ZVFrKCtdxHw
OX0VjGj2/qHWHspOITZHsOAPVVJC+/FK2QtQjy70aoTGQaKVQdElrB4oyHY30aO2
Jwn/grAV/pVl5w3ZJyLhR3ykC/pNmKxakzayywSzRSy27J+SN5+6gIvMikNKGgIk
UTCV4odlfUCKmcYJKR22s4hwNU8Knzpxn5gzmhahGtMH8cCJrjqYQXMgk2Gw4jCe
iKxfkgvPmUeje4OWjnO+Lq3qyxlIPhR9YiE7mRvtgRHPntBIwmPSMWXH2PrWdURf
g1hv34cHLosWwZJ5XXbtYJ1YarPyH8fxghO86sXLv6W8f7RTYplbFQpGp6Bn13Vx
WVCboIl3W63OqZ7Os9g6kBSa/AWvqTKvDdBLXA///suWxLQIqQKoLlbuU4qyz014
e3On+i3hTk9aJADGRLrUA63cYmR61pHdELbjAYfnrASMPWGNdGxoyJgUHuIU7KAt
7CieJeLmH2e5nZXXbxoWX5g04qdEZXyhD4whgFKM8CtIAhVCPFbhetP5suWUSgVL
PbaeAEoFb/vo206huzoidIO8Z/J/D/zqJKsffeSfuMUMgTUBRKO7+cXE9uzpzB8w
dqHz0xAlh6OQUb7PmkRP2yUj1EaAnN3cwgUMRPpDr3+NLni3ycfaF1DMjfqamvOM
CfKJhaA9l32P7OrYKEsnHDtJ1l78ixhv9jXaBXZDXWxICiJ32zavMrnk1YtvuE1R
SrQ6hyf/F1izRRez2iljwAgWO8ofDKRX1Zax+YxS0PtxrOlcgkJJ8k/2A0DOGk1E
tWX8H6wNtrqYkWaV714nqEEtG/ivO7QxI++eRqHEt1GdmKu41X2QVH7dO46b4/bD
pV8hgXLlsgweyesTyECj1zkYFYnDq1IqwH4dSqkuJWO1JUmBgrJ9ZSUP5/VEBkl7
81ljETIF626OrCaRQ5UY3qu6ZZc2J6bw/omjY9YuJkxhIIiD8iqPArhTJU9HQG0u
iwVLhe+hi/kYTe0ZBLyHASjeLK03+jsuFUUd+i4a3ul2MkDRmw5p9QDQBdQMxsza
wzb3b9iJARPxJmXdg9NZGefw75Vd55gwA3zh7lpTQ81MrM4qRM1ublMTPRXoavXR
POCefveIoyuiZTep5l6ZsVQz6tvAvY/MTlt+KILy8rAWRr8sH0u1Iit1GUoAdcCG
sJ5P+Q5IWSNEv1i9HB77tEIDI2hCTY/XrvmtyIFpCZKBux2tzYL44HlS2FHG9zU3
qPBL0wYaJkbkc4D2EDkpybDIzpupWc5oxiMDN3uD/g3DmpvkhhPVhF2Lc7FB5O9E
jsQKm7CJk8ZRUVslHbvfvXRFSU1eRuQ6fhoTVA2/FLD8zME1+IvGfjsXu9m+708r
ztEGF9Z16KnNo2ob/4smX+UGRKTYhWzuMJY4uSmIxN6pl/rZ7q9KtrfN/L+efzc/
j/ejQ0duVIee/GUjdDsV5u/MwCGoq4VAxP04n4jLnZLHPzX+Nn458AgadNzfX1gG
/6V8Yb6dbHS7ew44YGblpoBdZ3ComplsnlKfUAtXsz6R4urzShTSIKtN7YkZPPzy
EDiZG6unH4xPZc52fvzT9lVDAaCjGT8m2fUKmT4VHi9xiaDGwYelwjdslq2S90Az
or5xKeQa1si27ZPxqynrJvCYYAyfFTfQRpGdYYiXTnAwdIj216ZCufXV1iY555JH
bF/1r2Jxue7hhPOaLXzKmWgbEOKaj8aGVK1/4FNFuFLiSnsrhLgNOzcVYO/l7qDP
M0ENx/iyEcFzP8qIu785aXVlDXnYvYGMxaJLDXiWqbRW6prKazj8lEwM6gWnHvvS
YORJFE5yqpL67xcgAYopbRyDmA6yLk+LUTORBg//yzy0QBvFRhQeDtpD9RzgU6b+
KUEO71q69O451xiM0FAM8W5JlHb3s+MySrpRRN7ZC7/QZHcEAEvLAExSkVZF8TPc
oQ2M828FZ5uA80j942kRy+teecr1hPRNjAFG3EsGqTRN55FR4EXak6tzonrc2n+L
XKSmW0mZKFblZy7GkWfsYmA3a1sJ8D/fKysGRszG7r6foA22e6Ak1INClMdcn/oK
QifZdxpbyKcZQ6zP1QWEWJqutV+rN3z/vzfAV24nDkEN/mHqLMpRiIZFmrck3yTq
QLdhyiI6vXyyLjPd1XE4g1JMZImmWGi0+CUTGgoD7eW0btiwj7J8qip881bU3msS
w3uVswd9EaaP77dhjdIhXIsot4Tz80qWbxHYvaxFDo5MTcf9b71ABf1Bm2QJUlk6
0cl9kN9vuhwwDEEoGynWAoU0ImPHoF/sFdfrKGgIeFqQAW+3r07ZkKWoltRcc4eA
xx3E8nryuyskVLY7ao9g9X4sis6m6YHUABnVbjh7WZOEGjdRlgDjX5xeVBdSVFFc
FPcrLm+uXpmI3EkOqukWrgjVoOXXehuWEwOjb3F9NlHc3aJsulLbTLxlKdUUVZEn
GEq2VEIJvPIgwBwlaYNCee18OQEB5pNQv7Sz524NdDx89L0FMWp0/PSAKi1+LSnP
VZ/ocjoDTpIGS0Aexvm9LK4j+MPYj1tFr4GdTJFQUE9QcceUuuUhhjcpCwWmNfPh
xkEjDFO2onfs+gAl6WOuIyVb3EwOnaWbkfg0z0ReL1tssWE/epndAIP9S3hheP2G
VTc+45xQ1Oq44kPfBP4YzOgGcJrvTjDr9ZExBHmXXngKvepSiQ8G1bW12tgu85Ju
9BV5yyPiILeT4kslwnUu1NAAMLGh8jkPUr0mJ9Oq1TLwt1N84H7OYkmaHx7V9qUQ
inr68oU3gKhlj3Lii0LrKkh0qz03wEWl2uzxcz6lAGacEzlehyX/AGuZwXgwtLhz
+ZfhzMepTYfj40ZAEjXqUTbPmsHmmPEQh9LeOiHqgr5K1OW1TId5Grln/nHWzYvL
Au8p7TA2pGqm2jfCz2XkDw41cDmvsbLBOcIpqrXE7QXMc6N+Lsz7uFxfpeDkvjze
sT1mJTrP8SjA1IvdX1c1n76BcXcdwXwy1imC9yqw/QpAqAv5Xw1xriJlV0GwZpXI
lzl0gZoUvAtr8LtUkpe1xjwqMRunDgNVYGF+ZVhRMghWTJDlVMbbZGkIlUZDzpql
ljTIRICqRuYLI3NDqI5sEuB76yh88HT6m6vVMqZ9v0MrMSVMDLvnXEOeMTcy79Yk
U3NBaWu0YnWcjrGNDUmIaAo0HhCOt+NxdmmFH35Top4P25/QUwXzmqD4myg9kBNf
Vclv0XL80oF4v5XLiOE8dt6wX/7Ui+gZgMIp61UdVc4rZAfWwNNngmavpziLkwbe
Jzl7yyCxamNMYY9OLBmh1CJkY8qMoJe/uXMuAFqX+XuG0J1/mNpaHxfNgx9IsY73
S7ndppgSTZimQdLBn3JsTYZuyGiqw0sAwUAjcrGBCb+dx7FeHywaXqEAR6DJEoKx
3iVmFN7gUUUmt2N35ZOTClG6WEmUyXskum+uLlPVJ++LzfLDv0jmF4osXOfIgzvr
QmaBLEccDv8rPlu19SCyQt2f1tH6ezsqtBC+if8IMKerIrPPBjCFQAeX5yuUQjBj
QAgIADu+TPOe4ROgqBaxyvzAl+NHIRcPEb1iovu1TUUcMpFvuoemGH+S3pkPPfq+
I54VZpnoELzYOChj2OSq/7zIX3pa+M3R0usovReRTTeQTYk6gacLjBJnG8ZiIFf6
Sk6NYTJosUw3ilaZ9P6txkpwsGrrkRuxSt59HBf2r7gij72vjneBXRDBod183267
mr7O1jnTGpdyxk/9fOdB4uayObc1p9JLlSaJayBD3alHspsEcjsrixhkTuClnxBZ
faZd4xaKamsgM9s8gXGBengFUt8DlCpYHgwYWjzncFv/JXXMrn4YZXxiX1cRPM/b
R37ByjG9/oCj6G3P50vZmDY+MzR71DCFuS2Yzlz2+Ua/SMpWZ6sqqPlTRjLe+7JE
58Fa/5bw1EcXHEsVk1epANqHrXGUq/eY9K1DID7Hr2bOkpFfW0M2j2nOPvyc3VfR
0H+Wv2QhaXXjIGTdMoDWo4TibtTQf4INOwWsiSBA5Orw6//s4EsnQDx1IxMIhYoh
a4fbbtk+0i+7C4G3YhCc+wa23yxQxhPbM/+oSP0yfd8SH2K/04ftxK8VsXsbzEtk
m3EkdyR7tU18bCwt7L1ixwHIT10pgTxK/qAjLXRq099UrluD71BLJo+1yHdZmuol
ZI9CsebXFMW2zCePvsFUwmDDItO20qi1PJ6lvgPHKb8PeHKFB5X11FJSuytPJj6R
tdw9kx0WWb+yrh+jAvn0rJrtwRNyetJVvinU7xJvKxGn3aJPrFKhS3RZsnKg31Bh
gmnEMr12jel5IQTsYRva66XEGvX1bsE6RUrzrlyox9pvAoDTOZxmyUFBVVEvho35
qYLF5OOhRiH0dlD5YdPhlHBi3rSE+EDcRZ83e5E8q2kIksON+Y6KU+Lizr0sETWx
4Ojb+Y/DycHrKGbTfj5BGsSD8D0esrOtIFG7t8G+NjxmrMdakzN3mIlY6Dylc7nX
0BsQm+k8lnTiRYC4Ewjr4TXfZXY+PT1ifDixDOgIDFb3+/YRIMOYQHXrc9Rc64Ej
VPXPgklHxFMAOTdE5DivG9MArzPyy7PU23g/q+twzbrnjMAjT7q/H+8GA+wgIM76
BfxfUiY9z24Ec3YQlr1ahJI3tvYUK8A5JBo+pGD7CksAeH6PZ01SY1Gcbk36Shl1
dKutGks/TqNtaTPacjlzk4is4ptFLvdrpqWZWl2OBWD8ovJ9NufMTQjFL6qEBPaG
vWyzQVr+D7nPYtPW2tculwoBOreT/aOnG5aKzeNCWub+mgFE063IdZGV4rfSY315
e54pX0Ntz33fsFRaU8HZT3A39logr1soztZni/ZUFRYzVeQQ2JLVCW1iIdr83jN1
H9s6smW9Ylkft6Zwudwl724Onclyje9sJJg9FC6dRGd8K07KUfUqg1YHP+ZW1NtT
6aVyYa/qM8FMFOgN1ZcBP8BmGhnjLBx1upMY+OVno1aHnaM2lFXylzEYj0db+RZS
gVFaLE3gPrc5ZyB7vBEjP6nGqpom/orwfmFTbQPLJw7ooHUUAdvSeMLVrA8rYOkc
CbVjM8KkxTRn3IIfJOQKa3JlU1fZP8zuMCyrsH+eyIVcr+EZPtKYVxikItkJYBgW
cwwd3t9+a2nzLRb4pytcceuRnGF9jTJQpdPM1oE1zRsz1aMIE83ikabk5j/WafLT
GPjrUwg1MBHOWHQhjQ1pVSMNPhqeEGEv/Keho1bw3pasGUQV89aqA85eMzfwYCWH
AACvd8gEn+oTk7fMr/4Xx5y/F73VbDbzkxpYq7EQqXjUX7Kz7m30xQJ4NXfQM0PB
K3eoJrKFT8XpjWE8kI1loEPGnmWcUU9JFhrDTCicRENRrBuzI2fMqqPuxm0g21sW
M+YrU6Ajfug2Byu9bxtBsBOAnX5wvJPZa3rOZTnhH31YlIV5ji+7bT9nRGlZWG07
b3iflgwkHO6EoOyIEE2gwVSWAqb9kf7JrggGCsSPWCWy79MuOEZamwXFjyXmHvHQ
eJqNlLbOLAxHfVTN6PX24UyPq8Xf6i3hvGPKHyavI62B1KMy5XngFacLfzxoG1dV
Xlp0I7rTjCMJWkP2Y02+k37l+Hl+zumXC+6ZrYRPO6f9H6+Rh1GGSf1JCt+zxjec
uv6OIpjspjes6fkmh4gammhOjuexgAl5ZHxFCMC0OcWn5eMC6bowtdDKtU7d8Fzy
ZesSXiDhwinNGNqMyPYGBFDfu0MkqP92QNbkk6ReXRRhMiPkFxXuaPbWxLHx0css
uABnL1TcdBK0hs0dgYt86S7m+8WQSOO8dP+D+zp/ws5giLE6S+PMYgvsWzGI3+7+
w0MhHWkCyTBTItRR4AhI7Qt8om362bonYU+m/s3ivuHIR2DzT3sMDkwzJLx98Kz5
CcUYz97dqT34yMenJzRuVc46Oqg3igFu5fYmkDcMX0lkCxEbjgRsWXHVmZPKpcqm
wd/lB+NgMgUDsjfv3EPUPt4iYd8iBrLjkBY2b4z/T1UIzv0rNwBRUWyd+/NZefT6
xFE8Dqv6osjt1njq1TCmdc+2Qqta470587DDFIwlImHgPk97OoripCT4Rxj1h8pn
rx35m9CQo14994R142Hf4LsoaJMneC9mvwFfDPLCFPb7oGuM5A8hgz0Dgwa50uqj
uGHDjwXbMxm7h+ilEgosR/F8lhq1FGJCUa2sQ/DrC2qq4BWAXHKsy6ql/4RRiNxi
CY2Zlx5ViD6w81LxHVaA+o8DJt/enyLcKzYeaYm+3+FSmARwyp1yidtZmZxQs4C3
44JS72TNAmX2lWjht10YJwKVKwqJk2uZbUeKZgiV8QR9Q3s4QiQS6R+7XXc5friL
SXc0pziMp0hVK2naqJzJbxiB7wayPPlzk4B2BqnzidGQn+PX/Z5KX82sI2Yylq92
W2hX+oS6HOf6libWixfyAxDj9O0F3AVYJSIT239yUNOae24Zgo7rpYo3nj5+Mw+g
bwcukoCKO/0rkTMLdhSqdgLnss/gJAuBZ2cOkwQJP7kgC6wrpLpqi7Zhv06p6DZT
XRRQEN4eFckLMgx1fr5JWtrtXCnGx/X36vho+gRtqInOj7AV1fRjPLbqNfxK3FCV
vpjwDueF1ivqAUU5kUkSSqGm2n7l9JGwFxm89JT/xq5MJJHfmSLezyIHISnCybv2
d1KldhYLS2XAwlBVPljFSjLK5xAkcgXzaKJtd6YIA1o1BjKgYPG6yxLzh0DcqAtm
7Rk7sLdFuCX//O7G06/txwncj92LHaIcD+bHC/s6AuTb6kt4/bhPgbfbUic9rFrQ
WGo2KOZ75XUQw76h/0Qz2mxJOJFBjWhKtrMtCyunOTizo4noiCMOINy43KHnCVal
T4+9y3RZKT4gLp8dd6peOGu1tpUtoJxq0TMa0VcunSckeXGIcShEbcBTonQ00ayk
8ubvin/y62ogbVEIKiHWK9aC1NvXpRPCTd178U3CB8sZL4sTamMnFVyzBWpQGE+/
81C29PghjljmeszwaKZ5op0yb4nQIJCkqDxwgOJLQ6MGwu/Qmqq4GnEVdE4/whzO
Vj5U1JLu1RPfM0KF9PzmSIPK6Vq8HUQqinBei9CXq8n0PXKmO1L2DNqabpf8tmCS
y4q2GOmDS2x3yMRd7ZbWSE+PmGM+SA34PHc9vT3woobwrw0OPOHsE7sxPuR4aaR0
B7D5CgG2OrDHDwmxC3hQPbZFFEHuZnXHpiwlHfCc41NLzVKLdDHFEPGr3NyV9/eW
36Y/P/CbdKClD5hEdykrkSmxJ9MkmSXQ41VdQjLgnpipoF18PHYDllxyEkFKRy1y
PKKNM9ewWAhlnuHw7SXNBe7basUeyIaAEmZh1gGPfn88vJ+oTHUZBxKRRknKZGuG
35rc9q50pXmAkMMG0SqB49Tn96WwXvbXt9VOr7a1Cuh1GoantubliGjf3aK0LCmM
JkSku9v4nzZVbiy8oE67C2a94oBxHwvI3Va60BEKcbgEdlFNR6pICydky3QXy0BH
+hoQakFDhoWfN0GH9337HocsgjxffkLf3Vc1cYaNt012KVaDXobgGYV6URC0ZJmu
rSGOm8ac9cJuNZxza5RLPpTv8CZek+yQrPqz3yClu5iKopLSO7TmxJPMk19OTeO7
mftZKuehliEBDeqQ2fcrpfPb7qTHckDJ8gb1KgqFAhvkO/rs9Bkv8U0eJJyZ65kS
I/hwm6fp94EqOrqmLA4cZpvSu+t7vWHb7pSXhJhERG66aR/sN6sEYeFBVvt9pmWG
99qMYz5CFYap7iV0Pz58SlwysMyNepffS1cBebgqzzlc4KKXVem3HZG6SuV/YgJF
Rz6hy/Fpz+8vj8Pvv7rSXS5r78kQXbaihnWQvG52o6ZjbhTZ6cRoRmSsTFcosBeM
qiC9XUt7zqRykmqIEX7J8Thl4IXMZeWSfI0uVA5mp2SbOo3Cfpm/bjR75WTBEHEY
7o6eaIZRRMxvebfR4QG6Vt2gzLymL29EI+6j36qaqgTICimoLrTPnBIeoGaxSgBe
gLjVFGyHX5HxVzMG1YqI71X7yLLfFfcQ6+9A3SRUfcLR8+GcTsFMGMgp4nAW0XT9
j6LqCsX2d9isEz0hAUAfGCPQw+PlO0h9jEgA6s+3nLrzx4oSf/fwH4w/aUxZ35Qu
4utHHeK77S8+v51eXUgbFUCGn23n+tTBqrWKm0BOmC2KgXVsWnpU0nkm/Z9v/HgK
eJEroVWVCQ65xJqtGPm8uDA2FJLDDbcWIjo12nvaw/KIOx7LxHCsR5v+yMGFRz+F
MIcyPknKVC0Tvccdki2qJaMkyq7tz5wbWXtcc/oYN19a0QiB+hgy8rtHRppmM0kd
kfc5B7ZPsurqBIzVEyzlyU1434r/xpZK4CTfyf1w9zhMhf7IvjYfT0LyIhOVC8VZ
qwiSufPrXfxOCW1vKKB0vxZup+KxQDyn489G2t5EEfv23KKLVjzajyY5NTiay//C
4kAbZFr/A04dEwFzYG5jjYORXSSfyRlss7llv/HA0PVkmxz9FHe7ZA4KAxRNSxEg
RIpSdlKDOkHf8pqe8rdJB3CEnqA1PzeHLavS6bTWsxeojrZmWmenNdMhjJKro/of
4IshpoGoCe+MkRS7zPhWrjBIOrhOTaV+ARu25uD5o05LGnP0jLyqxX2IH0e5P7Zq
roHWPrxveM/KHOLiRYbz7GAQmnrMhDtOkIB2Cgg5ZgJBe8XofH5xmfz7ZF4AhztI
7Ktdrnbs2Ikq3HqFLBVj4RjGbcw4+EysXtYMSnnxkGcU5G6T6NkkEMGBQxn49rP7
D5KjizyrnFCNGFOPpWegNmYJUZcQtRhIUJTj9E2wocarLyDuiNc4hNWoFdanfeVf
aTE+lYyivOvKDVEkTHwOF5ONB4zeJsaBSF61JxupJbf0FRtpRje1QDb5RxBdX/5R
KTX80xL7MFOCu1lF5/t2fU/35IcdH9NeQhVNGC6BUX0XRDheuF20xGMugrFXkVYA
D4KTuEdthYQ89zi7NtZ4WHKND6ehlKkcyoY81T97mX2PpC0HH4P9e6KDJhIBZQpT
uyOdR3LMSCu20CrkqPqLw2EMymmLjUdJ+H33Jc8y6qjczN4dV6TMU2ngdVuRgscM
1nVN7Ojoa7bi8jktNmKvk0jvAIpaiTTImZILcJCdMgs/Sqenj7jZtFxCOnNob0I+
us106AxfKsnvS7Msuf351jcVRmH6Bi9sJ6i504SCh2N91m94lUw4G3hk0paCnEDM
Ggl8PCG+Pb16GUB8vv5zoRgWfPkJwVlRURyPnNdDebNRTlEouDqfbA+PCVGmlvsi
XOGYSNly8YdiQHsOpVLGrw2TYCoKzAmYNMBziPzl1aZKvYKGMtRm9Zs/j8LV8bjz
bmQ0r7U8wI0rphd+wKHATJEVSoLU+pQJFFNU/l4oC2f+esAVhwfw2tSNwKdRAhFN
NRdW7lzkkGR+8UIk8L8R8m/hRedEMn2vldOR81k+96PIIllNqPbdaZm5YJnzRssd
t0c0VIzpfMy0rmHWFb6jqoeSScm0B4lS8w0ppbEPVeFgtxsUYq9LKcLsfQl1mWKx
/M4QJEzANsGkbdMDiXBz8TYGxjsiFXXdJkkPDi7THrYqFGLniKBgMJ/0Ul02Ay6X
SlpUATCVyCcLzrRADEU9L6jcL1y5Qt8E3xMfURL4emFuUz4zJciEh/eBS6+6oWbu
wqjnouL/1ymUQMStQxzygOkt0shXXsADDF6xLmGcTYrd4AFCxYpTyQlUmBNsGNpy
441btaAZhNs2T8dz3FplzCAyQCRbxgpNaMv6hkSe+611exRgZVWSmxbzgC2VRqrx
bJ5I9pHxRjymvn0UMvA5POxBHSjvHvOss8rAJ2R5GAozWWM5ee37ZevUq1+I7bsi
cfRVlZOMNQoEl+Wdh2a+PHL9NqQUoDAkPrvzlXXPgmrRy2SY0H7YjKLlVbdYinyn
co7FuoldTSNzOveAlX2nWWaNzf70vwmrnA3yvrop43EYC8M5LuatIUh75hW0khsZ
aWMZFHPPzucxKpt+M7fULwAfusJE/86mioBn37Hjtmt83LraeVBo4TWRBlCvsn6i
IW9Twu62mrZ8h47qOYK+bJCnwetR1jkoJ4pjn37HGwzcwgYqnlmCtZ5Gr5ng1oDg
suVcY1RjV1XckB6t++kuzvbf4odv6VANKu8gEakhHu6fJFWqpTXjlLm0KQu1FTtk
bRln+3ZZBN6S3ylTg6632kdeclY8Lz4hSrZ9Ez0eSvVxbODvnXMbzrE7Jf7/J8WE
iXiwCAHzvVffqfr8FRD1SAnWa6mxrxiQEc8o7tekPdBQSFtlH1kyIt/yrUnAG6of
7JKPbL6lTSMfBhrTCzYITvRMzesKcua76hApRmgDfkuQav4JvXNoezBV1zp1VCeF
siqh6KPLvmjsjqCYpqZqogJiIHePjQvTg4gKD+kMVHvO95esbOp8GvocidG+em2J
RQ9qSmcxa8bsHqDsUYyr3qOOC995UVxDPZxXJd5C2EcPRhov6G7QclMrtrC1KlnK
Pl8i0xkX8ne5YKzv8MJpmWlmZE8UeHfDBtCjBO5FKoOckxiOm1QE3gnzLxH4/IKA
6l4+6tnWWPB4zmOBI+8ieVO6WwVjA9Ll3pfEwwTGP3taJMaXlJQT1HWMRfm9JoY0
+i58ifi8/L2j9O7Ut4ib0iEEWzWQfZ7c1M9paq7hqtzKsrb8V9JEBPTJuL9hkqEs
DEzEx7o/XKXdhVNErE2vQTj/9bbX4XnFc0Yx+hjav3fI9ssiiyfQgPVhTmOzkp3N
/DWpiNJlMi6e0y4/0PhL7uB/56qDE0SYL//ZL681r3WCpYzq5IPbpnDwh6qs89lS
7ILEQnH1bT3mZFZG7hkewouFW3YFvdreCl7kYIb6Pp3A0YRdeHkPfxQ0AmmTL0kT
mgaqWQyDhWDVyIKLx8KRRsoz/K6r75pNqO21+zwhsubW+SzNKH+qIycxPpz/khsl
6fgMd8FLEQGOucmQbrSc9WUSk7BlAxf+HtyQfDk0+2tm5q1KMfdnG4mJXT6e6GBi
1ge4HLDBL7F7ugZ/w3uGcEGHm4x0+VyFTYZQVHODi1ReZarubm7n0mMGswEDTkXJ
W2TQLztMi5JfBDNADEJ4j9UoKWA+4+s5f7P/3S4I07emxHXe4dTg8k/cKQOJgJoD
jokvVLmQNFMJzyHwiSFfUyVVX4n1CSL97427iS3Z/7XsD2WPGvCv8JGag61jV3mX
x5QRt6DYsmm9olhsEJqHez0MF92NsOaF0CWsMIHXOmHNoi9Fa2CKZ46SSP0CBoWI
AOSanNh7Gi1+AJOSCl2qN2SrQBYso2Nuv0i2tb2pWl6TV31OAM5Gbdy0YzGKrMF0
h/Vm82s6JoPH+OGX/IXqBDVfIAa5ooxd4Zbpg66xwadP+YkxSp4vXkMA8t9nPDHQ
KWSAUt6cI7ZzCvXNYGBkounhf2QAV8TWobytzPE02aNNdWzFzz7E6V7lYGb+TMF1
bJtuPlaxIz51BYrpVWvNhlVSyTJ6vSijpJ5DlIzd9cybuXsgbjVGtEImJXuN/l/M
5pWnpIn88xDsjkZ6Kkt/TeOxgMA27UniarEzuQzRfF0XDAbsdnPfLxK764VemHAD
Z+x5D3cWvQaj1sAdAXv13QKjsDPugIfdV+D8ENoAf2u0g5946USa3f0nt3GB5IBj
X+Sj0CNXbJcTnECYC48MwTW9N1lMoJ1Ei3tElv9SzlPXnJyPoUOeK/MycVuI5Cpp
xDBn7uvAzNZRKCiO89cOImP6OdZ5MovrbugajF1KPFcgNy7pP/r0gMaPORggzx0t
6Y+1EAv3ke0Wyjzu/XG6cCyZ4P4i1KbtAHYFZl/e/rIRwLnuFUzVKQnAaA9haOc7
KpHl5vhsOq7tUKtqEIoiw1qnomBMniMFx/5jwJhoP/aCnKn/nnrjvNJnk3NZc3UP
5ql3q4WaHKgH0NgGBHr5FoWWA80dL7EtJGRyA2I6f9wC+BIFFkRFK4IIqrkFfo58
85RxRmmPCowIey8UqiTqjzvd7Py2jeWESTkO+fZ2wCEsdkZSy2h5J89pHbmBS7un
`pragma protect end_protected
