// (C) 2001-2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
b6CkvAlwkNI/9qTWdONhTf1PyBgJKdrBrqY2T+kRDtk7i0cjTw1d3Qz05UpqYKJXLxwuxfbWf4He
2Z5ZqD6/6F1ANoJiECnVU+pgKeuJ9Jh3V8KGhHvN3bgV4qMofiHs9cKOjMdk/dH+amTdHQyWualF
45JK7f1FBcV87CCSG4nXWcPEiPL7LwOQ5kwnTROyPAxUgk918ETTZ7wbP/m/eD+uViIbTFlEYS2o
RVnnphBHb6zbUyRAclmIXeAoUOH87ArcONuuNB2BDrMf4a5NRYp6ng7gNNo1KdZmMNA7LZ47yguQ
HX+6nIkZJWew/xDTl/iw5jNksrO/hTWGSL6mQQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5760)
zwlsUsS9bexvCKMdanTiFy57TxDwezm6kZwjOLCopZ2g7tiDjg3MF0AiBJlWc7fNBbZ6NIBPBQ1l
wDUqQVoBrtA1e+Gpmakbz1p+pz5dqKxSWXVRslia3/bstz4KgjPNBw8mhzOV4XUqp1wxmNnqyMaz
XvXHQ4Xgnh+uMW1Ntrx3ladCOMAFEo5AyvJSKbV68qz88zVDLPyd2cmS21iNdV4IlO4CqOVkSXRG
KksQP5/1pJhiGDMgcgvR8hD3TmWfJKO85PFAo7G1TtW41sKCYvJ0vO0r95uzyV63JSr04hO6wupN
WnqpRKhKvcwWlXDLFaqajL+ou+A8dDDwtvS1HzWn4q++NMru+lvdguJ5hPoxRRyoUdTiJ6e3DGcH
Mjka/4ywmBMMD4+gU8h5xIz+ooM9BHVSHlRTsNh1orukYQo2UColP6r6Hs8l7PjvkVriBC3AAu+b
T7JDZzXmBStPU2x9HbXWaOADaT1KzdXyC8p+WD3qQtBJouM1QqR0lz7kEcecYNrMp52awC1ezKhg
THHPRG+X+Wft42ZzM9nXQXnmeCp03hDo21workzxThWxxNcO7c+qYQXTWeSwaiDChdwIp9D22Owm
yoBMtFXXpLeQuOLIpiO1MmcqnySPLqUt+AC3tk/EyrEBPUhjBfN+qOb+XWV22JJif3kLs3Vlnfn2
pHFScAqGuGhAnT0m412NQtP++9HZgWY1ibLVQMU+wMv5gT8buK8I7mFLzkZjJTSLHsyhD60rR7ic
D5ARdm9KyFcCAP2Y4oP8/4HfHLlLqSc28UxA/3+/pM0d+EhXKKGNEHTkCWzUto1inzVr9shU4XnF
OcR7B+NvC/tHZdgif4kXRd9Qsx/xZbAxsTToVITMeainPfg9ONytiYPi9VXpVDEcGYP/cAvfkW31
U6DrCGWDq8x17victTyuvamcCPsDGXgLfDAn2Bfjmohu4nIfH+GSmar/+wd3/QdvtWCgZq1TQ3Us
XC/6hi0qvTtqUvYkCCVRuCeA8LyVq6tsNL94P33OFN6+/M/VyNwWFJdcEJrlCKupJ5cQi7A8Sqnv
uJmpViB+VznFwauLVWPa8tQXUrRvj+SbukGALYvpWNHMQhJdjbv1vQ6vsE4oiXuIrNx1p55kr/xH
xzIskDGOBXEZhyF2B/HCc8JPoE7m8qoGLI9DcQDphlFNjDVXtzva5XttSw5fna5hVXpxsTSpY6Io
Sov6SNkhalMBTHNdpy1eD/Efevw/zpBesYdrJ/Kw/GTLiRr/K4b4iXFqiriDBjsz8h118e2JKN8D
ZpEIJVUSiQuFrPdyYxq2yr2zzojyndSsRgiHJZUZjbiuxMSzbf2bg+OpDvek5YLw6UoBuJ/XKyfX
3fuTgwGHr6jqcw+z/EU/Do3GZihjq6S0TEKtTysck5aO6YmKYKCSM5V8gX1vGgVxyIExklnzZdqY
4uLpMZSSQIErscoxH3CKtkPFRDjbpHtD4NXe/VxIIYze+I9GX76z5QtAzSeUvKC0iet525WAhGnK
wD6eiHMyAXQqYMCMDUhrwVrKk+91Otc0myshWphn8NW3TVY/m45LYr4oncNn6EAw08eKEmrl8Ka2
TzCPvy25McNgYdmMu7PZFLj7UTrwXO5yizTAeZrbKPpQAmaNIY/JkmXecT60OgJhslXA94q9MeUu
Eg8DpjTV0M6O5D2qMdWL6CqBAiAkFBZenRjEs1SDwJf0cDtQwKtBU8VqP68pngBm4/Ohqg56ku9K
HTx82gHpbuoNQSJP0KddR7GTYqbOFq8Y33IRaiik8nYWOJ8RMFxY0nISuNE3pTBFt7w6e1wtOH8e
asA3jlbbW9X/0T4lVI+fP4WxvUAMtpdFz5/RZia6zxUeIyQSF80C5BSXOX9hZpLSnuM4bX/rAfZn
b/O9lQI+vuyCMBf3SUnUy9po5FnWftfUkuHJrkFSAiorIKoA0WOjAYGGVgYTUjMkOZFi1MRZla+U
JQ++HE5bCaocJ+JDvOPXZ9K2SJibfJoOmOfaoIH0dM5gznWnWhmAWrKYPV4C19dUO5tLJUbEl77S
JL+2YZc7zSAeP4SGDh+3i9PFQ91zeZFnbqA/Agnwnk3tanNpXAJbQdBpluLmNbhDwiWxRGC2mfta
j3MxHafwm/W+QM0xLjNM4o01W9tCIAXsRlUwbuCTNkV8+D53vOIJEOFOmf50+zZslwy1x8sXL24V
XDEjbDshaYR0A8eS0wBhRwK5hKwe9AWuPo46oLluVA9qQ0RR/nCLGGM5rmDxdaZ2f7gCSbcRaQTA
EUPdQaI3O4JcqM0tQhYqFKkRJcIdECAEtkfZBnUjwIPEAK4PY7tLS7fa+isOdwSWNrUF1n9Kxfb7
qnC2R7fjifUPdoz9SJMro6ip2W3xeqJUmbgE1myUOYgHR05Myi8YPJO1Ck+JMWr09+jXHjslLTIs
B4kReShb9dlJue/rFlKwfREojyRSENeMOEXKMDfIL9IJIFAGWfZRpTcJOlYksARL34d7BSZSOMXY
PEN8BOtMpOnZvSo0mHIKQww9fiAtjVwK37qMBS4McVbvS8TrLL4emdohOmdrLLeHtbrALgYP/Nbk
rRXEL+tJqJS//dX0dkdrl6YkkIIROCODccGbenZRIOk7vrAS5rg/7l2v2c8EIZGrHmfexK4OPIxm
0+4kBA+nbb/R6trBWT3CUWFkPBQS11MeRTqy31r3uWW2HkOquagEggSfEitFrtMETonWk4YVdqJE
ih5A4o0FYKiFe+x18fC1nj4O+kdPbrW6f3VmKelmL2Kjz8UrZc4NlUhIfFMr3vewrBOQQjV7BTpZ
EonhfzIFhgc5v2FUs2Ox/UE4sT6hkXvlAnpCgp2S1N8m4Xpd97dIOujYIamA3+IrgayjkXiM0rLM
pjtdVFHiFpgwGmgv5GX/+tv0tvUGZqdVdQRaVH/KOnT9Q6wr9SYhmrk7A4K20IjjBaqQm9z8l2mF
zcGgc7o/J/XcClxGbsXuI0ZfRS0NxAuKpSWSCKg+RQXzp0lVK+FJipXJRVF//spk9WlqedMIp7Tp
LsuSlIXp2i3ymk+39G2z1YR5R0tYbrzWr7oc8dcZUmcLvgKOfyAwC8Oh3Rct3I8292JiEj1gzOCl
bCA8fcoTbixi1pR6F6w6TXpnnB5yV+ctrR6Gk9t7ValPKjQAIW8/WA1HZLmnS0YVrpCWT8nCuM70
czbBxphfHO26K/4r10fwaUZIEhlQ75WXdyYEQR4XZzVPBH/ewu0MINqi5yccvxDdKt30OsQaD/Qm
7psR7TV+AI0WDlmGIzQjIUbX/OsBZB1DYDqRU0up7J4t6pvZgWLDRDWi9DXuMPJ/kLsAdKQKGbSM
66g5by2BCBSOS2tUKXmiaF4mnOKXnwxt+swFjGDpt3B5CIUtnxKt+eTCr6utxyPuHWRMss9I5DXi
uWcrevSAaLgYb4zvmVPsmk7Qkbzz/SoFNgDD1LpkNOuIfJWsF8tRO/FBc7g5P6qaWwoUjLo21QYs
ubctOccyhGCS9omiMF+uySthxAZFR79JoX0AmAI9EYAqPJ4xWzgd3xdZuROxPlmI7LNjrI6dxFt5
1GPc/TReuHPLkdB4w4m7yE34dtw3fPt3ngEcE9XM+SrAWuKIB3strKaiSBN3jPwDIsKnuUUg71Cl
nxHvRxt7BxewwEcGCQD8DlwAtPUmWtklTzxmO4RQQRLKuOSBiZJTBfOu5vascTTCeYrbNBw0Sx8q
eE0vU7rrDcdQh1AKwwSWhVoZa2XbEd7vyF9IxAhQZYiUt/DzGSk+GswkDSrICB65/HsaYVYll/53
Ht2Or9nf4/woM+wqGNIcFe+kgNgHgZDAP/Chc/aRBIikS3p6fGFy1YYPCcWg7hsuPDLtQdol0eUy
Q0tDfbS3zX+ifxGytA5xSf2I7haByBW2wYDn2mRo/mHBatgX5uSyPm06cx6h7flCxspjp9sjGqqF
Oh9AWUJ9ALhsXyQxhGiFhDff8A/O45P2cvhr53Kj5JZBYNKVCUUPCSOHVm4uABUfta3oIfNigGKB
Aegp2sq1OX7QvZnGE40racyR7D7HrcxnQL9nXULs7CqoQuXUj4sfLHwT6VTpnozeKy4WovgYcRbI
xzTyvhHnEHap0jvxESE+NiIb1bouvxI4RfPvMrrUsBCg1++bgFqAsRSg3x7X5bhBa3E5KuNUi3cD
GGZ7tbvrdQ6NAViQGpQsOHDGcxzHrVM2X5y1TNEfi5zc1I7ecZf8Xs6Ebo4ivJ+aYAnm7QNB2Gi4
CEyvOo4u6OjcD3dL7EeUgGYBt1jUPiMhehQooKVhNDYAR3ISb+ltahM2T68yxp6/TSO/BXHbURWQ
5+sXo977369XdqvlpuxCyVus/6rKixQArjaS26QL5bKTMUirMzWaf9w1vFtWVpyxhl7A+aRfdTY3
BpHunKrvPLgFVYK7Lrj9oI6pJh3uzu8jODZSiEZXzEyKxlbvj2rAjMceYHwGgTMDMGI2zFm8oKrj
hOKo2XB177rlcOKttAK0KT8fwhZDf2ymER6JTStYKUhfOovJNRniU1GR+FEGlAYkR6ue7LehF3Ta
epLemtf+5Yq1pJhoUrb4YQzdrIhsAdsffAgon+cphLsWyREQEW7lJplIRyyQcmlrVcpN7fiFw8G3
FLiqpARwkCbn548EI1Zfvo4aPEjbCHY1Rq9wMmFYgZdOlTzUfPRpg07iUZRS4Aiwku/yOI1b3Djt
IRkLC+IdEYIY50ZuDXLDmujawzOWjjbXrJCWtRwCzaC2V90PEhjFc4eQeQh0R9/5LH/BkQ20OxBS
ad/LfF/Znq2yjoughu3x0X3rKJ2BmdM5oTnfphIr391jnA/JDl0PVBV9sI9m0jYNctRqkMoGQiHr
InRvC3JxBFDRLN8b5WUD43NQJUITPqX3Pk0EdS9lXXmqZNpLQS5i2J76jhyWrb4x1/qXyCaoz3k/
vMI0INQ5p5jy5vsL0PCEC+ALiQp5s0J02IbqelVy3A2ARjVAPqRLuyBORdmDiZNnyKq0E3pXiOWI
XWbhouOkd4oDnvPArqKbzS2omGvzWOHPNmAF8baocnGP9gOmbhVXpBOvkZ7KoFl4iKmoW9+K6R2o
G8Eios+Zo8gu1PT+Ox+EL5KpOLpCxR8qMI3i+2as/+aNWD58zJNQSFPRY6cRwVdkrvLxkHAeDEyi
bfBygoH8aEAQ2T/9cAFGXBD+1kMem3cAC8Ao9O53cvdjJmbBhm8xEZwvmCkIQlIi+l0zBVGwt5HT
khV0zpmi3kz3iGFFxnMwD3Pz2z6pMN/tPmwe/ngUUp/YVA9gqi7UhEU2UEUnxLb6ooKIhIQR8iNB
sF1fEf91cdKcsxyt+7ehyxK3mxtj+VIGWN0myzREV9tH1DYZxfv7BbEc9yOldOHFMbMIWeMlyH0y
Q6WPOsjNzIGHn4U0XH5juQBJJPciYjW6OQkOiyEzGK94SsPrQwpauBYaIw076mAjAJY2r7zCaT1v
1cmeOPJKRvmESKW6wZ0xuMgWUU4u6Wshj11xfMCatVyc9fUk7xbl8R8GQ0SRGHBLCMUDs3wH8foX
lBImepTty4rHnH0gthiWv9kDplIrq5Sxq1oQsGH6iWoxBM9OGEJu4MjaC+Phmodva7U1zdTAfoGE
XuT4NANlkynQNntMZcKmibVjdyqSC+vyxo+ZLYA7diCgtiYM81hObmR5G0vUnunrMlwUYEFHQgxG
xMhQjoIcNqwlzpga2pta72uXqmH2VUFnmHwnjA7LZj5qjmiSKjWEH7Y1agNNJXSXU/4o6tJUcP2Q
kk92wEgViGLK6By1b+eghWKK+IBbhFEvTTUkym9Ora3XOKWyBIr7m8k0e0EokjFHWSD59Ua4V7D5
6Cl7WC1cIwp9YpBS/8eafTX7eXUUhmMtyWoYmh5gsPsYyyQBgCtZAtiCNo94emGfUnf07THtybrK
x3as8uj46s2byYwZI+iPE7XdHohZKxvmMDLrDOPUwT4WF3NPfCnF9HmIDyKZz/sa9mHUoj6VRyry
qUM2siT191WQ2N5O1zL/npsxOvCZ4q5Hd0zVCr+PkUrNjFH7M/hF2R+ohwL662uwTXOfr19oduP4
4R7PjEefD6xZVnBGUAx1Y+VcBaWEPZTppUR0gJawoTgNqAf5X3xp+hpNSPQLmVTCQ61QW3EcyP+d
MDK9V7uQO2pU6g2E2wAx6VoEefUv51d5qBkOXpfnZn01DoDh78/vjSC7xZbHHSAVaom0qm75mtg7
DbUc9pdPDlaVb/6SZ8XaZbYomsmAH6hVx6maqii6xny9qdFlWFy4lAscxLg8lqZepnKzqyr0fy6s
NCIqTsyXg0foBiv4aman/O8xxe8y5wdZ4dp3HW/evbsKA6YiTUnZDkOO79xTmQQeZIdrwA6oCTSQ
IYvuE8ruwZCEREQkWlMFix6NT0/IRwFnpNbHm2YI5LcrNWhqa2YaosOLJ0h+uPMmBwJ/WKjvTAjl
ONUVIO6MnR1nPKrZg551giIyo/abJcTRo4V4hTAvQqJ+HqCLoRci10nadBF5fK5Shalol0Rqrj41
FqJe3nMmR8RZzjbFI1wYCR9cJjnR1CnkZZKdtUdxIs2j8HJCor9AM5p5eoMVD6f8NilxekwEZLTw
SaNzXakqtKdJO+9OIdotygbAWmu5FG2tRRc2imHDXINjEjGkvWNgw3KLzZ64q31zrSh+zWeZPck3
KHDwNh9Hz7Cfa+WY9CxFK30/x8UnIQebcAJBAN7zAargY/vjvyVZ+Vqup0WHS0DwLmhu1b+7bApS
/cC+GyZGakYRjQdlJo4ll80mK3v2U4h10ZblEYQ2u5Q6mvFCvGgExqOZcjGObDzZufOFyqLbm8iA
M893kB7BFMa+fdKb3j8F8PABNHXX1nZP7h7JkJTeNPEW+hVNslg2tnWNxODXsCGudRlzCPB+TE4K
wdozz7LdrZ297g64cI3ulRfCEQhJxY/Z0gP47xJzvj1olBDYlqfQIXC5B0bw/JKffFLv+oNGn/qf
hB7IYbU+6RtR6MTciAgFBvNdaYaE98aRJXKZz7ns5ZPYQsMqsQQKCMKWhf2dA6LiMV5rV+1vYrzr
Ndz6xv0M8K98uYWWmV8Z9UQDGBNCfHUrfFDg42VqCpqFwAZZWld3P8QEeW3VeuSUXZV2Dc55uXWP
Iu/jpM06F/rLFFQwd+N41nhDtycYTRdA1ep6mLGLrR4T9H38a6xAazLTNVAwEDAbm5aixfhyBVxW
WsT/0UpMFGneteyW/Smu+vP4L/4gRr9rNvsjluKG3chGYQTZNnzU4eg7jMsWDW8nmeWC3JD7DSds
Q6xM7Ydcr6texcaBJixmE0GYdsVlPJmHEq+DgT5GTTmCgnjTWZhHC9KmK1YIioHDoPxNzewGnxfx
epL83WB+25KJ0C0rObZo6PvRDts5sYaZ9RvQea4K3+NcarbTP/RoOlc89Munxja2OfU3L5F+YXws
EJLwX7vdSGE3liB+Zl27ftzdALzw5ZiB3SzeoXPeZvBDFQxmRp2oFXBQkKozFIkBwjPI2r8zyZGs
kSZb7y/sHDErY0Y0RP5Ry6BYvWMnro7uaxSfj4M+H8wHl6ZZ+padY+IsZPv1SB2bTFN5lwvAiB5E
LO104hRjs3Hd/ujqBiVlFzLLWlZnREOHKQJ5AICSkoqJNMoL6ZwNzVxWf0DrKwZO9/y/ccUCS205
pQs3
`pragma protect end_protected
