// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
mIiZPDkqKsoXS3POSXEwVBwKxwpAe/ypG7UFwwM54DM0yncFSTQsUqfFat5C9r493hPin2AmKdgB
BbVlsyIZP2KSFn3H5qfmw4I8EUO3NAPZlRdfJfcwNlgLqWM5dyMcjiogrEzQW6tuzZo2QfbBcsgP
GP5PDFSv2SLNziZqATpGpIjBFrc4T8mQWi8ZDAOBlyaFgUS2VLT1jr/mldlZUvzNkMX129PtDAnR
j3OrLgc1qMyN3F7/xRCNRVK2BkN9POnF8hkwic0f4iL3xC5gZeBtHAubXzKKIYgBmJy9bOQKz9mf
517eF55z4yTAmeoQJLCFm+9+qGItqSwh9tbQnA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
KQJa2R1thyR9CzK7NF2fkkRvhR3rY1V9o97/KTbzxgat5WTQo/vd4lNmGYNh4QHn+J8hU2k+3XsF
iCsMrdT2gwhpQQU8LYl9EeOGxIaMU40m9ugiHKfYLI3+12SAfrwTCwtbUh/gwGO6mMQz++aeH94Y
OVxWnVz4J84mHFjyqpKDY58vPNW+SiKd0wjmfRbGaD83g9N0iYJwLqYHmN3gvosboisB+yK+IFy/
UZ47D3Q7eovbUu3mrJcJyzQ6mj8lCnaZ+K5nEXgOh8xs16UtQ15KKHTLNUlUABHG4tBXkxdenKS5
rtgHLvJkqdpzZwrTSedM3SMvTOK58sUSST586naP3HlgppRiVh+S4ViWxuOibOn5IqVGWgE/0wLc
9mmEpVIQ5vPMxAyytBbe0QyiyVpRGohgSYYLFo7ZjR3sp6wL6dHqgZYAD2fiToMtrTJCZpJH2EHi
b7e65Kw5azVJceO5GuFMb/ke61rOHz+9DnEofz1+Mx7feiidWwkXu6ZXOjipvdZBr/lUvaz3h5bw
JA572ytbrvLvlgy/96mG1wCO9LmfvcjMBZyvtC6tR0wTZhKQ65bteIoQB8iSiUwtwP6LqQmfXnv1
yVKst7lElkrMBFudAXW+7Ncexl7Nb9CTlpboV1jCm7FAcDg3prvfshJatoMrcsh1WRpumzhB5EJu
BvBvsl20hjkUdI0/GCF1E1N5hrYsIw9kVTc6q++shlKYvCtxjYtSsNs3Us//z2ZTAK1fl7YWebMq
mOcvtfznb73Mu5SAEBM80n6lMGE1qDyMBjjhwZsmJXNjTyhtQRly9MBGZvMgRyOzJjzLrWwAI8LI
3TxHGvM+YtmLBBYr6toTvOC7skCO8rIJLB/tt2na0iPDhfen7LV18LIySw4NrJakHDphLsOzcrnf
rCIx3BEmz9f8ZOWW8QlFnRyQ25Lu5D9j1KV0k+XZjnCpknxOp+++wD/+tooYpG2N/DIYJn3hg+Nx
Ud4gU5VcACjlrN1I/fa7mhb/RCILu7SxQ9O6M/OpFs0ylc4YwpcwLLX38Fa+rS9zm940eedsigR6
N5LYdUSo8kpkdGKEg0OlNFyi3V+b4uT+bly7Gkt8/ij9DodWOD9P4XQQ3GDae0LaACWQ5eNb+hyZ
LD1opmQCaGWNW2N63ErgNV86la6O1BLmdilxmfOVbASmCrorGPlBBHQFX0e1qJKsUpyOOQxwSW3b
ATjeu8QTg8NnYIlxPpg4CAAlQH57EuTuP9yR8igDYkyfa9CMEIJu7QC7lfTB6BmKUEw1YzkjPpS7
a1NzIQyedjhx0tcnti1CdBDLlSnyXXjlHqRjq27tVeQVHw90QP0kRErFyrJLts00l070emSCBGUD
m0wdfPal2SZdi1eWPQYimFUWx88PEAmjLfSzyjy0HJQUrlHqqo8qAR2f/rQ7hACZkE08FfZM8j/k
5Du+c0NX6qfQrYCQgStrTD/9qJRONGaqTckL5ZjVFGuhKnmkJcKaRu/kSwKI8zITJ7NCztMj83K+
qMGimFvqs1xcyATw8XQie9rNhnV5e4NS/6fNL4okHQ6KqhPeE55cjNRbWCoJtN2Sh3xEmzbbLuBb
7nDfP0Zf/ms3AtCLVzu25P3j2NzXXOT0WDwgE7XO4wHVrS0dOVsogqmf8bllAoWImopQLcbZsh/s
Xvcq2AzVc8R+npDuLjRpeNnv7ABfr7fX+zRW9ToN2gXnohXI/Ml9ji5gQ3KQnm4zPC2hkJ8GnxUy
zU656Q2hm+uCUrt3Kvd7PyOBoEgPowamEC3vRyyRlBtQKsui0lYT8gfLOdLAcC5GF+NhbaQw+fGa
MZIO5DvE+290SdAoBYOX/pmD4yJ8WlPvHV6Z6RijfV29fWuG7th3raQClleWQfHCoUau+d5vsSzA
AfaCXE5bv2dp01zbKksjW4fdunSd0cYQ8CXlLAT0g2eaXbH+bDpRqMb7J66qlhWG0l/P4JiCm8n5
ldoK8yRrOfALc8Q8uSt84ud4s0NqaMAcYRbA6jPQf52GiNPpVYrzdWXf6Zygg/BxT9ZGBjL47g0U
zVHuPv/JZv4VmGvAGp/eM48eUYSpQlneS2fj/ieLjc8Ha39FeNf5ObwoVwtHCe1wvMw+u3UkqNtS
1cLBlaSXOWyMz7dwD9NMMdA1HniS6Mlkqssbj5j2l/FHleZMUhhY0mNe2IunnHGy6Lq7bEso3Vfk
8VdzCro86bC74ySmZWtU4QOaWJXXAcM/0SPr/YWCji+m4hNur+lO67Noz4zDo1HDiH8lx2Thm+V8
ucfWoximaQXe7YAIyOniFrB1I3NhBCLS281+ERNy7cNq77bfkeyUgVAdyoEuzDX9GjmZoYH5b0L8
LzyfilbAMdJkhTL6MsVS4+FqHqAAFdVBLmsw7jCWjzWlZeyPI0oZAl1enK9mWhmacI6aWXtJInMv
aPSqyFOWA0XKmGAB2VVabi9dDSAqQ2NgnVryNqrn5IVKm/6oB6snY6hIvQ7WAqvh7RyCcj5trvCQ
sGejY4qGMymIdpludgzcJMy/jh1X33vHXAyJtHKSR5G8wD2cBUAdL0gkWsf9lHDyIngm2MODLDVg
McyuXMpwCixp0kXh4f0eSI9Na0GkJ7kwmo2PJzt7mDsujDflLlA+L+NQn34P14UoiXEZpKuu/V5V
nZPsBsnOxi8vagOu/Mi3/4r0msNp2r1C+sh6dxmok0Ddn1T3kWGbl/CIBaH6z6nX+Qx8SVuVt2y/
28rhV4Nl70B/+G9PHuMoNiEE1lj5nXDMzNTsYE3pfrp3Zmal2w9bIVPLV93BdXey/M+ba9j2v2q/
bs38hsy3siVtGYFgnA+BdFI8I12Vi6Vbdxmo1FPCrYzjZaXlZbk6KW2sHfB88ggceueV23w8zfRI
z+g99GShIokdZBMo1S2R1k/mhiOduzHHksVl6hw8gyG3AItRrbmUcLfza4QITJoenAZ1Av4Kbo8/
Alkn5KRCr76UgnRrYYmG4lHN3R1BdzczYLiBGMxZIkPFfPLOiHc0zSJEp46ANXPSbpZC2uGJs6ST
2D6dEf0P0QrA0XYgujq9km98Z4Xdv+5EiwrH3Acc3My2ZgPqHw6K5nUH5gN3ZCAYJxQNL/joLzGD
2OcKXCoV7DdXmHf1duxELdpd8qdKEamGO07BkUDOld8hElJZ6zhxVuEunUHi11aBz8XwozeJc/BT
SNI2ugUaPZzuiTiqX+jH/CZ4qoSpVYoZQI98zSFw3vs81RGjtfYwEmHOaBWv0j2ZDq4p/ApmvCSn
oWdFkknxnVkq3ZI2rp2Pyg226HjEVGou8Gg5v9MkucwkjI6ESdxCJ03n48inQlB/cNy8AjFQXGxH
BA900A5i5EAQMGNrNb6mMQRwsi57GEQP9FAEWhp50XK9c+VI2/FsbzWTRPD8L7NeNklVTm/E1dsL
1eZpJyQ5PzN28sWh+heuOWatnHgof8GFBCVmpgAxG3aAsXz6fY8gDbCbiukz7bFYpzfHZgo9OBEf
o14zSY99KZY0ziDmMxnfHznWRIBbyIDyiluUMuL+qo+HMBtHcw2bg8FLSd10bcCIk3VcCWmAihkr
M/CFinlhQ2OfVOYtZnDKRLH10j9za8xYyvbX5vsm6/Ohqd+R7Zg7lbpJvH23dMcKuAvgadiDQkEh
uNGWUWTniOoDMDiWTIdo1/4S9UE49c21dzWmvjZgA/CiuxLhIrIMeTAus4FfSgu5xzt+11/dPxRy
GnPlI1sLepnYVAUTcHldpydlZfjV+XyPjnbQf/KKSCfJH+bwnjV/EXVSGYOZnOm+5vmdWW620YwO
QVpYbOde+bVyxb2QpOhX5VbkqzaNnVSZ84C1ykifgV/+iIg2nDYBcNIiAIO80THOljz+ynj3y7jV
wbd5mOjZB+y8kcP8Kg7HMUb+OuPE0c9HYBSPZQlJPEHbGADveetqz5zxTwzxD3LKQ7e2zKq3tDHr
WcjKQL8Oui3jJ4TDQOVgu/nYzrZRtBcdRsbcCa4KdYKOpv3wm6yhhJza9dlqJNZHDoRZOyM24K8j
sGz8bzxBFDpYgHKMBCvBjfEKffE8Ft37WLB+n4JHxIYDAs7ccdFTsW2vYFF6frZeWw5qYGvw0Po+
L7KyrDkan9r5A8u7VhbbtkelUvSMl2oY/XIadIMrEAglLL2JhCxQoVGVizGRvdcIUYYUK2tVL7u7
Prw5a8cHnjx2ZECdiN9KxZ2xnfehj9tzy2Zb2Q0IPf8H/J/fMEwYu26TujovVpgddh1G3n4pIgeR
goP998Bygnsz0z+M3jq17CJx6oYw31ilm0C+2+i9LR8aJT/jed7g6N7kDi21u0IV5niRBMvrM3ld
GrtdCQJeKUOva7uTHdaSVzYyr9aJ56tyK1ljPQqvZQvUKRsRJpxiUhwRNu1QLjUU/+snXoG8gBYT
KNxBc3+5HPApf6EUAnxH+Wmd+QL1kgMvpD9NyLeSj8paRSzrLfM1/VmyWo/tXGdjI/uCXN6zsTX3
/GykI27vz2U6jbL7A48JTQ5qjvNV+hr7g0tG7Bh1EDLANoTPcCCXfwvEwYBh0xkBSm+0SaArRYA1
Ckgbn8VfR5MDWwM1PxAujDSQBJ0Oy1SyjR3wFQykvG8AR0ffTPPOdPpq3r13ZhzFXhACcQwex5Fe
y4Ga/xe5HrOlxwCBIP314hWZbdR2MxdldWsDmEQ+dJkh/KZ7UVZPeQwHu21uJfN6S055NAv7hntU
PHy0cOK4ecfgREmzF3VxAks+TkdvVlBMcbYvlMt6fEPQ6iqxe/F1FFF0Ky+hjl5avuzSeqWM2Qp3
6/wJGBHFdI/jtTuRgVCT+OM/T4DsP1f6nosxfgo+33StK8QIHyi9mxhY8U7aFs5/nlb07uFSYFCg
rxRihm0JShfxaNjg/p+TgkHOrwZgNmjUVtKPJuO1zsD+C+V9SZEPUn73BYBzX36GphmLWa3bUn//
oB6RXpd+GPyaiwz6mxnyc+4NjOqoK9eo34q27+jHnAbf8HcFy01o1c9lfQg5mmeKVtW6hFZjVy2N
w5bmJx4XpLQJDArq1yGZV9oQEeyFy9CSV34yzy299GvV2QY9Oke+inmDVYFsxlp8uAfOFu+WLGa8
rFd35uQyhzTu38fiHlyEXY+7QGuqqg7W7VCp47ApHVFx1QEyLL5eEy64qVWfKhO0juQgCClmBbsj
mxIhGAO+cROSrVhuoY7lZyvtq24D9dv/SjVIKzEPho6k+nIEo7I/NEioms33GLUN55BnbwsTqT6+
YhMDJs7T+xplpAit1riuH5iHxpDOxv/Pp5RXil9deRq3lYzF+0VE9yCBj2bBT/Zy24zppPW27gRq
AxylL/vTpOSqYKzjNXgJfO5m6KoFg8SrbOlBsCVz5+/jOMHBkB/6RCrGFY6SRpYmSmu0xzuRqquD
fOzIoJ74h0zdJwZLulhK4sPas1GfYXDn3CpVvVolyQGuypPEcRmbPB10TwZV7Wq/tIhviZS3sYW+
+oq4ODrnBeMOPdp0ti6yqO6FMu5xS3FPLb5pxJWqkndJUN1DlfI55RQuTOeRmWrvXqoM/ntIS6l5
ViHYtqmwNBLrLRvi6Yu7rZIK7boJAwzZ9/wVjf42JLE49hlNCB56e0OPZkVGnEg5MxBCGjtKoKBA
0C894/3FgCW2+CkyaOOQtqdCPO5q1YO1AXQhJ2n+ukfrNKxPVWxEKUIElXSqt5K0wJ5KzCjnQddC
VGjUCzT09B49gQC80aSYsrGbqJ4I/nT4x7NyWQ+hs7MzAW1jBbfMOwqRPw5V64RR+D/GKKTtFWsi
fvocgC4ECeguLi3antXDhp0Pak6sWPvUTTJNy44Kyk0itbfnp1AamUaWJYKCkPqh+MzF8FrwIic+
+kfaM809xeU5jeDgKo0vl2wVZmegsckaRlISTL/e2B4ih045/VYSV0EK1CEy+vdm69N/JL5cRaSz
iVrgDwe1yix5G2Wzq5l2HOhHpyZqw5c6cjsP267H79ogtl2X5vk3Ee91aHrseI+Zr0LcRPKQv2jY
SMgzQyjUOcb33ql+yq2I3IUlfJZemmbaoqHkYYWfgjK7M1XJEgo4IwvA+47TEx+1F7HJra6Z2Jes
IMHtK9N19MZr0HmbFJ2uUzQo+fY2VWVgYK1oUz5+CgcD39/V/vbARg6WGPmkUQr4Zt1AjUawfC/8
aMiniiZAThunEbfSEdJ41J8Oa7bYMQKT5OEP5TNSfhS6uvfadhAu/pGzdnzTz8gyd41yQb3yPWPV
jTStFsSVtXoS4zc76SaHfZ5t4cE+GRfGsf7TxggTCofwt+jLh1XQR5MBcjfG4eGl6aflIu6vQUXq
Shxg4WxNMkFXXUmFIRr/ufNAeADc92OP9Zoqzcr52GVwaUVBQoXZ2MkKrl0Avq3FPNXIgwf6eb/e
fCHNHm7x36iceZMNH2YwJMIFarJVwGpU25WHaDjX2jEb7YBl9AgQFrDf8F7/8o5sJjDwpF2KmDNA
2nVmZ6bL0JwgJs+SeYoWqd218ZonETNjF9SJtzBX2wEqtQiFnlgBmc9iHIxg7DLXuLU13+t/2b2Q
BqhLD0IlFVPHclEHAhXSJFNheYIHegILbyLUGVevJU55Cx4DpFHhhKd6/dGCJK7Fnj/Q8fLvyrdO
V9cMo/z100gVLUMQ6CRdsso//ij1MizBq6Smd/WXZ66Z7G0BXR5CxnzOVS7I4QnjO8Lx+L021mlo
Exqe9SZ+WBjAfq6Yy2gIbbgFs+zi/AJ6C7qaKjm9Zo6WitK740vR3B9Ajpp6K4hLxx0HgXrjKoh5
g0EUvkkpde/v809gscZC4bhHdPU3aciRjKJc2EtulhdwjTGhGeBvjqrLNzZ6dO2nq74DuukbV0Tq
tgQ7IUHnKbKlJtPHYNCykv4HRG9hwf19K/wI1A+k1mYv8UTfgutiD0a/3whX1MfPzYMV2LkDzvxG
Yepv4z3jT30oZqqV80/nrhj0YnI/gfA7eSlbK8bzaMsfeWO1DQ+UgeAnpgBZNOmKwDVLHcEDkwE4
rF9srWPxaJB2nAFheBXG8Zl8ha8=
`pragma protect end_protected
