// Copyright (C) 1991-2014 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1.4
// ALTERA_TIMESTAMP:Thu Mar 13 15:23:43 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lw5w9f7dR7Y1XgaHIUM3yF8yag+eDxd9MRXJqIO5PD3S5VWWcHXXPNUQg+NOUOey
hkdlOKEKRMGzcrzHXlJqw1Y/03zAH/OGo2XE0RGLKozXVTV2FdKWh9IUwcRTcvx4
dkGAPwFCykVD/Vc4j0fQKLJWk+LY9hRC1lRf9u0fk5o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11264)
CEKQjQlKC6CiWyTm7+IvtezY4t39Nb+eai28Bvi7HsjGcmpJcbavetuv9US2RlaY
mpcBxQF+VqpfdAD2cqm6/HPJaLt5HRUjbKMiLQtnjw/5dCLAFyzBR7bDuEb4n9UH
DR0Y8n+TgrM8znM9C9Dli91XAtvLZWl9zSW6Kjx6EIwsE+EX692dAXFULytWptrw
TyIWHqu8WFaJIKamvtDZ+9EqdRlbmWlgf/U0k2zrekCHjw/O68Mmz9jREmrmaZHe
A9TjYXIsb7ZV92Js7/NA7nysSCFpW070PTf0EscP577YoHbbPkh4ue0Nk7qCvGIA
qnKu2c4AVMp0X+Mb2cgBOqID7oOFjdN8RrQnc/YyFnKwq3X51sj4Lud9fMf2DizF
GQYCySR/HUuWuc6RaxdrI+1tfJZugRXrtW74JYU1ANa8JkoYgFzwkwk6Sx273aXO
nhZb9Vt1lhuC0t1f1rr3fpafQO9fwDmv9L6Ex922Il8bXyammMo77LAbuWPgroWj
zNoAB/qaBApkO3mpY8aDwHLAy1+mMG6eA85bJduyLKX9vqPO6MhRZIKfRumhmrG4
QlkwWzddmyx9c1x16NfEb2KUvsuCtQWrsq/KnCfuH4xvQmZj0Tfo2cWhWOOQXvY/
pmDHMKf79JUFS/TzFL49NHDTKl9Xj4eLLFtv2zZ25sVfG2/9wt+75KNVHNsAADyn
2UgyVxuUfXCrUji/oIBB/xxBxsqofVzfOXlEdjX01IEdb8vX2Y7/B8HOZ2J+eifD
VCRn+6COy3SnfncN42I8CpedXAVbq8+3pRIZmZ6RyUtezhf8KIzCmSr5ksCTPdiY
zkTWTjcLhsEs5tTyV7urGg/Eq/6WsUGqr3ZuZWxwN1Nj0thudAjwji6VrUT/mXyC
FuiGH1wTn2HzSFoqhDkgh4aX8u3k+mhrt+VlECoq3jBMbLjrjg472I9uP5yB8s3z
7VqeC1rSPRc6zNeNMPWmiLrLPqfOGds+lyu0ZRY3R3CMPBgJesXO2E2p6vH5Cj1A
Q0ia7dUYA3eSfVDEXr0Cw8PY9boLcbk9nedppIgvMnt9if1ZVjHcrOYd+XkvKd1S
F/DSQ5k5af5lvKbmHkqFuRJtNCeJQQk0x0WERg11svZqk/xTpoluC2GKsZOifyyQ
lpf/WkjBY/ulRP2eiEoEGCL6uVlYBiiLwh000ytNpdOiN9ReREBL1Rrby42Jpl7S
vLHSmmu0fneen54wqK2b7ymqwuQvAhYmefG6GOVEbyQbxzUm7tC2XGDZVa/WGp9/
tt0VDWTmaqak+zI04HauZ6CPIhDFna9v2H52mV+eJl9HFfTFRV2kV5Tqqcs22I3M
W+kwXH271+u5HxTRKIVJdU1FqwR7fgVvQDYsmezAgZJQfcmoUXfTqPMbHfC4mgNM
d+7iDFrCyEpaXob+VFdSOOdilbkiOD7qccR5GYpSLHVgHLS/dD92D8BTijyEnJqH
AGmtUmjgSz8FsmE8tNLNQs/Hda0lffJc6T4DqjbYbIxJd7nCt7j9LXfR9iIprNNy
liStwcrXiJXWYXSCuk+oSopMjY+6HV8bnHMHpF9b5oglFpWAZHzjXmibs9dgA3xI
oduRROyNZw7lJ4FMdYcXJEf/kDCP+eCa1VFe/8gkn9D7DeCw4616+0Gn1kPOllJA
lxUxY3y0JH8Xpor56bC51BE7MknqD2jY0tC0sBSIauM2Rl+Z1hamuwfrNrrnYCkd
6u2RLA3X60krelyIC5X8C2dW7kRRoC6iZhxRUwuMoZf2Ohu9wULS34EhrCGsbax2
2nFE9miFTP93Bz8s+573aZGPB0jeFRTqG3tALaGSKWS+1EeO5/U0p9bK0c7iZagJ
2djdWizNGdIVx6Z5vy7AZiqqMPmBJSkhpWsn8fLennsUTVt00U7En7ze/iX5tul9
o3kCvAGLsvI113qNZIPLtQ0ktKLgjzK/jtJHQgO1cCGqhTo4Ro3pPVn3LhEpDoeR
ibW4LEpt1HMd0aeffzUfFeM4eBHQPcbpwxdNpwAC1hdE98BQol14HUb23RpABG+R
CabKhz63//VcXSSSuGovPPc28RQ5OlY5dccSSiJhDUo3t844DUZzPkniP68Vty34
oMov9t9U48AY+uVb77nhQy0lM/R2ZxMJFkRVP9LknPf4KGXj8DPlGu+PKv1irNwL
9eESxzwKY6PkSarb3IPXh3sLb0WvTq7logYw5zhfICkVLJuOxJOm6AuHP58iixwS
uM7NnBysZx2KYtWkaECjjXgyOBIRiXL2r8hy4BkSBlrT8fvIczxdq6T+o1FlnP56
n3klv3Lznzsncbs2fJAimht/yA/e9JulXSiOr1VsVg6pR8huBYo3TlGUymioSGRt
oEkrwCtFPB+b26588CNlJO5wYjUqp9+od4+ZgYSHxWukmUfBaU3068wf0NRxwaT5
24LR9bkaCkiyW9M/wvH+TJF+ASuhgkCXF5iwD8c6GCs2wiok735EMLZFgJssSGbs
I6ddZJSwqvd/icAuTHgDTKH26JnVKsSA64FVREbmAdWuU/IevlQeX2hE5NIXXi7x
gGgibiMrayy7LvFk0oO+jo9WmU66ltSDThefkOkQHkFTR3o1K4tlBjaJ991KvpCG
Q6ALvhrCjo0nKGWP3OcHga3BHC8SZVT0KUSLqaMB0dHozp/exAZ6/kv+FjbQmyur
20qDE3qIKUI2U3l8kN8o0utflAahqFXM/gafnlQuMN3rSdg1BTCCbcJ16coHD8/d
yMyC+LhVVTyCWzlJGPSYr4yB7AUFBNZhE2wy9rhdcmoqmCntxGu19ASO0Pf3oPQg
UZFRPLYb4VkO7W2m6EqBtIhcDw4sESCWNemk0WymWfJ9H5xViPQnypkqhCrr3gqB
oZ1Da6F79eBtxJZiOyElIf1nV1QkyyNvTgJfh34bhGihLF62ssIApA49gI1kHc4i
cJqxJtsKEsajAtT+3VyNdKYWBOREm9x57jfqj64IR30m4FSMrClOTli6ka5gA+0L
w8l/rLNTtMAL51bxZRRJda2Hz6D8MNE828ysa9Q4+vzRFRUTgHAV21aVDvv8urSf
5iQPVyLNRWzg/Tnnc1/niLmm5kIxMtPLceZLu0J35EAWZ0XMcyYlBUhHmmCsKGpi
Dzy4esAF0VPyaumbjlk/h6nIJowKG8aOFcWhbE2xk9JfabZCSnDcRw3qvKbfBbc9
IEFw3FqBZNOznwzh49TFgMVGXQQz+1mBBMPUeQCkghHnZLORYe6IZOXvrUHc7FSd
6mNtEzms8av1XEyxEQfo+yZv70Dum4dvyzk2HWEiU6mDHySvR0E97Nht+JTzwQBO
rko6lZwF5HwMA5ABYTf8bC3+TVc9LFkOprtbRDVUJHTNs+B2ZhEAtr4Gx2ZzrCc7
BWqlW9vjQTPAj62as39ZNP7pyJcQ1GbhAngSlzrE0WwEBc/C6ar/eavJixV1wcm8
yzxqb4c7GnoQT0S9CN7rZrG+s3SdFUUlrms4J/k2EdcDQUK02TENE18hqTqJtNr+
DKKziZExDAe6dXWukLFVn5fng5JAepafS0liq/G8xuyi/YBWAuE6i9DqnT5hHYCk
FOp8NalFQ1BgvzcH13Y51onrV9UZiyUwsmqIOiBu2m4Uy5vqbiiaGYINH927p/oC
6yjFD2t0wl+Pue5py0JPDca9KnmLBXHxd3a4md2hxhPgCNGBfT5/t+mD3Vqhfb1w
fP1Isg4IAmNyVdO8eX445rXCzBT6ItRawtxd+cFOdLu9dr80kwG1KYftSzuwC9oy
dNP/MSDPMzPMqUItgBF4BD9NM411F59cGiVWmACaVvZzH3vtAS62oi/HgOlAmUEQ
IGLgNHYqMN+guuSgOrLZIUXl2vhA/IwiG5lbGCEaFlNtE5HoC7mLB/jo3A9oA1Az
k03L5JExsDEf2OvGrK6WrxnCBKxa39c8lwmSt2yOufI3g6CZFxKyi51tWEmdGWH4
v0aw3c5Sd8intoX7iiG3YhP9HZ2Od/dpALqj5C70y6nhr7KmnL6taO1nwCAqWQWj
m7wlI/CBgTYkix424vzEEtgTu+7WY8cTb1t8jfI5Ew9Ux/Ro4zeq73qaWJ0GkonV
n8sEAgmctE0KSlXqRcJ8NVapTrKRx6UhGfXDfErl7ECK2x596oZlhAZUye29DHPu
TGy15M140uvd4q8RNuwCWQl2Ynq9WiJFGQSGt2iSf6krfYWOtE6OQoKj14/FzP0E
9bST3GbJA4dGuFColSq4GQxdfyONWlRmknvR6GgDkXf21IW1bBAwFRaZ6aBaHTCh
yqOu73TEtIqiqrCH9L3/0Ri3SOw4T0dFc6HktEtmDu7OGv0AcchbbMvcvlzGPG8i
oCt/wHq5QZL9eqr52b5cPSPQKQDZN5gvyEtT5W53+VxywtCC3Pkch+0YFDXGagMO
sGBcV9wBftwykf9mp8Xeg9Jyesodaw19q/5gVDCR07sT24kgarpkdQnJkln9E6Vw
MnvvFpotwRf+akZxG976oWeQa/1CpGPUVEp8hpWBPAHBeiShB3gowz4nmmlK+Cvm
2BppFq8jBmrVsKbXBRwSvyRXhAp2CcR7OU1O9VYQzctLoKdMDIZi06nPAl6b4diy
U5DU5m88X9XK6ZbiSsZ4bGQvypIyVSNEvhw5Up1QV7dafKylXFe9Mbvr2f5Sy9sf
m+3VpFX+Imzcn6ipAgpUhlXn+WKBDUxHkRqVh2gekchU6S8nmrRODtks050c/UG3
q4fMmx1sIPjy8yjBerGVY/jXg8/m7irG4C+e9TwkFjXOMALFRQk0Z3BggZ133bRA
nr4N8AzRXOlUP+qEy0tVwJn5yG3aHENTj9AnNhLfg5BIomJ+plIIccopX+qwcLNd
Mp7mGnFsaEcFKIhgyrgO2+6vCK/OyBq0es9q3cruYyr2rSG9/tcVJNRtHeOgnD7x
63c5ugCZ2xMXUmNCRclWXS16e5nXxnsAeEeB9OR8aI6qsTD6gg+fOQMD80+eTzWi
qwcMNLW7C5UmqpB/M9nSdiW5wmGPipx+P2eOtTL3/s4KcCjt5tVrW4rdu1KRYuS1
++kgsojeTSwze0I6SQVggPo6MvQ9E3ZqUWXctdAx5v0Ygxn+u25SMw5eLur5767R
zVl/WC046hstGS6Uu+YG8ClTBalPLffXWzE0lZpXF0sF2X31XaOZ+K+Xuyp+2Uxi
XDUZPbySx2610EHTYh3hocctmp8sxll6aLhmfcOUXf1HkNaRC6x99QKzcRXnGUda
zdnjKrSfHCChNVGSl5my9LyxBYbgjGMEwgLDGT9MbbDOvN3IG+r2cojn+eDT1LiE
kI1ZP6MlWgkejmp7ZMbfpY+CngQVUOUxeoEPPnbgx+NDY6paWd1MY08FgqCVkDxp
Cb2BivkndggZyo/LnDWrTr77Z07YvzaL5lQLQGf+gzGuYURk1DnMBypsXwEOpzOl
mewLHprENCW2WwYgiNmbwyjz3G5jiTGjPJSWOtOahKg2mH84SCavwgyEw9BQqYff
AVYOUtufv/zZ3ixsNbmylhWT2RCn7B1AVpGaPUTWnkEbUolodc7UhWKVAbpNE57u
eBQ5E3LtguCY0QnvGqjUgywEE0899r/DnRaNcEn8PwdkWB3wes5Kw8sovefdUrQM
x4XU7CU31aqBrhz1A2wT4mHe82HeOFYYOme2j0wfKij0EckgXS2cx5bDbW9hDTQ7
/13k68JZNvMejvWXJ4/pYIyEuDhMcBICB+dAPrwJHVFfMOrHRJljEsxRr0HJVxC7
QhAhyi7SbDpC0VZUZvoOD3aubS/OzObtY77qN/ptSGHpg9YxsykIJ9qbguHeXxnT
fQX/K8+2sbQDtdZO3Ey1tYDt9j+U7FcMMLXIhfdrn2dg+nJloh906rG8luKfKdQK
OP1uYZMDcfjQUjq68GhOoax+V0jSicNeReAnT6d6vJEtaqODX0LI9ocSuNztvoME
/AF9dPikE43E4JcjfYBF4nUaBg9uZbLhrDX3CSngcKl+ffL6uBryM+50dT8oeDOJ
x6OIMBGvMzD3zppWQCVhzeiBp+Cpu/toIuXEm+We6pw7r+37zAKzUI4axLGoCAWo
/oq9g/4rpE//bskiacAcscyrupvbSOTGIMQFXPQdlmMl2nwDD4xeW6cIZ3SZK5jv
Aq7CxtoDp2/XVpsh1oWK4qv7NI9RM1l3P3vShQP//z1LOzRiAFESSZ2bpQ5gp1HT
c/O8c27/i/uJ/X3DzNQKGe9016jylzL3JbjHTwRQFZpuumUpVCUJt06DCCDEnjvf
lRYPx8xbKrqhILCJEHdFGeAMyA15iipfF2VNMU7xd6U64ZLosVt0+JXBIlTsNvuJ
mK9rUlk2W4NmSX8GV+2dLkTY4rhr5r5/Vdp5m61sjYhqDiu287P/l4/QZo6nIVrF
vNZLasAgdfTFjH17uhMh8QleXjBrFaLF0EY5POCRbhYoZ1JsF6YBOMxS1uAkbibO
a1PKGw34xBUTQlt5XAvh6X3mWVOHk7FaZ31C+WrGun59BYIpnQF17gy/H8Xy19QI
KAQR9pUH9Fm5u51iKqPYxpqVMSvFkXddfKVoIUNoX4Bv7wAE+bZ7zKlkERpgRsbF
aSn/kGeMLRQ1qKfxurw3fIyv/mojZ3OqjkrtEkT+ExolQPzMngnzPY+sLvehk4P4
iORemRm1WboPMlm/Jiwqpoumvf18FHr264eUudxOKrUdxhRZVelbUIyn7ApEt043
+zucIcTvuCp7kdcnLMFq9KXQneMcZV94QKsqHUwXxGNl8gaZHnTDxi5Gq28T+7Xu
9MtXsmOcJki/cJquQbgTcOlKNTCJUzSMapD2j+a8JeoO/Cfnp/FFRc6cLsdHV0zt
5B6lYhIuJ48IqqUufQ8Xvdk//4drJ0wnb9lbMD1o6/pvy8fAOOzm/o7nUYmnqByU
mZdJ72NU+WFvtZa9xnhUa+LuO6ay5yJfHfhn93kQLXJR0nuUSyTdpdkQSkBdbrSK
J37aKUayarTiYZTwpeyvHVpzG0nnfb2cwJ5CzUuOPhPG2F0K2I7odTWJxFciKDe5
RPBfTj+Cd6eraYP1o3dana9fwqgEWgRzSDN/ekT7eZZHoVC/y9d+uKpJzjnKwS0m
W2YYToincZT7pYd+GM5nmfS6yztvUMk0hPBgbjL8sG9KSWpNozWITqlNO4dnFmxf
aGIFeWkraLKdHTO7sKHp6CoKwy2VaS9r5JN3tSHbJp56TKykBAjBRymEZm070HY6
6q6meNZxBSB7+gF3PAzBfGCjQt3JF0+IXgVRplRlCJNIf2Tp8g0yxMbP5Ae947dd
ckwRn+8+TVq4CYkubczcLDPVQLXfcD/TzKiGU0W6cnIZl2kitm/Hl4BKJLTqgM5h
1wIxML5wY4QeiB0QgalwFa7bEUVMYGWPDZqaJdhCa1a8G5pMF7/DmBCD7tcQkEYU
32JLCXn6Pt03NRwz9jH7nackqUMG7OcAPpxqjNfYzbKj1kS9CoAsfwSzHXHPY8k/
IsemztFarxBC9iDAc2Qk19nMx9vwoAz4a/L+xuyr7AsH1eFApZQPLBIUYsSohvud
YA0hqILpdu8RBSa6RsCQ4IIYdBeoXVDjhlCoxUAgEsAnYRUGybbyF5VCir/LycqA
th7TBxKohOzWFQfnw+IinCa7Rs4SWRBPNw8nTyvt9JOueNWurYa5pRme7mJpRThs
MOYtCJ0a9UfKiKG8slCFtdYOBu4C3a2P+caFGIQ3pF4QER8KlDZsBCaaTPzaQfR8
LgmgeOiJPmWRQYCskL7boSK3XC1vyhfIoQqepw1FVeT3LSE1PvnQcSWpjwpzM9cw
paNjZTFm4y0XSFnvXdL5ydZO5xD1msdCue25qJsSeHubwadLca/CCa8yrvZu8b6z
IZ6aIiBVXwZDlxEw76XuOPvR5yfcL/c5Q6M/qWuGuOAetAehFF49Nk8sLqiQzgYJ
+/9dXT6ZyiEIzTlEGO3JvcIf1woLu5bzphV4WwrnMDGDSDGJMD97QpX/7Ni6kXEQ
tNbPa6+tZ96OULOQRHhluy5BH714iRTpxjF3RFFt/WnjAB0Pcm0XOJN8eLt48Pmu
rEVhfE/y9/lNB4tlOUMMz3suJHAOo9T7TTEy7/snTaJPFbFtzoUfPoOtN7yNQ/8G
GzvVYYZJ++eh2qf5HJ71QaHV9wFu+lUsFceA9kF6v5f1Izryp8YSAW0UJ0CIP83s
p06zU0FhiuiwepDjruexJaa9d+MsDBObxAzD6PeKGJTl4Tw3d47hFAoKXjsxeLbY
0nHqFWRH+migwqMEcMUwvIGMr/sSVhwm2Z/i7nu/J1PLVZFll+IOMpBHDyFbQHrP
2bPYboHMcQ5FUXeQAbPoo4zKBs5sSJC9RvmHwbTPYsOWLoatetYU1RfJvjZGF1pj
kRsUCWGU9XZ8oL4hzrQwylIAu497c9GCEMEOn5xYyy4QEAGKE+1s8QxN44oJjcS8
hYR5u0C54b1Yb4k7YhggtkRaX26dSzB6fWVk3U7ASbLG0Wb9MX6jh136AvwlzfXJ
Y45H0j9o7US2qc/mlg6rW8OcxPLuDHc3Xa3q6gSS2/uUnmSWwOAgINzSNo/MRMif
X2gwRJaKVDXMGzPS/KFpZ6RtRMXjZmBXJvDAXR83BHMAQ0GhuT0Hrk41UFMkSaq/
vUgZaX3Hhcfz0xyy6mp+UBivG/9dzscuyezZFrJRqk55raKl2tgo2ncXRgvAU/sB
OcFRDeHjC3jWlD/KVp49nuEjo4MLGmF/4+MKtch3gXfY9eUexJyD30Y0MfhUCTJo
uVhAwIgLqyAkDbkEFD5X6cljA+GBba1ZmruupO6XF09XYC0ASJmw8PryUdjT187u
wHuWPOfsGFIqdMFuGoaRadQUP+xZawsN6tOWKCOZj/1nfqZ3//NZ4/v+UJ2t9fZP
MbjRBKs4BZS5lWFYs/kKCowcV0/Uc/ocda1VDVhT0pOWsNcvOeEuKFusdB8SWE0w
UhAMcdhHbn79MapEF4uYVslccvcDjsgYxBsbAA4GRaIW/8DhZHQ+DP7e0QCsoh1M
VS5T4QTW2JIsNvMr7nBR1LHnkn3GT8IYPeoJdgBQ+yE/MYMQ9nULCDM2+hUaLl+/
hv0RbVfZNCKPAwIaqxQ6yPJiFic/gKP65SC/FTXkK9f/FI8HpMEYxFjNg/aGLKjV
9jq4Y6Z2CDpbz6Zzv/aFlB15sbtU0ic3aeQUdenfVVlM4YyyOQmy0FLP24MoxECd
dKq7wDuGt9LmuM235ZQS+m2s7gubokEh0HwFgSJQKctwfJCMBFX0J4712RpajsKb
4WiObe39EwbeB4L9VvpT3BWRBzEhORqbJtdpYA6z/2eL/KFogjeVXxdNGJs0fp8/
sqkZnGXTJHEeneXlE0OOq8+1BC24iDKzzvsuVLloEz+Av1oUNYYHZcalXiymmQcn
oDXEh0HOA1CF6F+yILVQkQb8AzZ0VrIdH+2dbYw1t/YTdQ4pON/YGu9f+YYe2dLo
WeSfn1mULHwIAZQdYr8s+WRvb9HdjfmyNLZz8beQv5XJeAJE3SRJkNw0KeeLlXYb
r/yGJss4wpshqnOzzNG/fUooUGcW0+Xf//qzyIrnH5Dg5vjd7fzdVRNydn15HE9j
L8ShnYZ2MA3+AqQTN+DqX41gsZ+pmeSzTSY5ku3YeRLDcopebQ2BaT2h317Gnf+0
0TWLw3fEqaut7xxrN2QmIUb0k5vq6TqFEM7SB+LgCjdEXFOttf914Jt0lMtVNKco
T5tvCMqhmjI13IJcr6LyL4zIP7L9T9f+RPKdlUzdm25Sm6urAebE1rA5nme7HuO/
zCNC9sJgIrChfUwpBQEaK6kbB55OPv1EzAhjJB6mH4GiWLfzm51bS7bOReV/waVM
oPdO5nriH/HoDGVTrwNb5/9FfnB6Ex9F+/gVUbB/9PEiPujVX1WSDJMNTTYKccn2
S4uyXKcCPL7JU4KdRI8zZ4pvyqFaBHNMI+BY3vSSkc1/FU5Can8VJnR29Fvgy5VE
r3yrr6Y9JtgcCcbNzS3lQs2FdZDue/copvRkyC/iv4ImWD1I2/CTapyDuGkCAk72
c76ljQpxSb8THjBEdjn3aNcuVJYMV9E7SVO/ZB3QEFU8+BBu8XJkuFl62QUAY54f
9cmMkKTVtr71X4OTF0g6lEWT4jttbo3Ha2XWwwNk/ONr6QOJ659en/lwPLSihNLu
3uJjo6kT5egydtBVAkWyfhwQ9InDFdAoDZopjNNyNKujlO9iWpVATEDvkd+uMPSh
YWrOZXLbyVor2JbA+a9WaplgAqXU8Wj2yYou5dkwgoi9CNd1OQYRlzltt/8Sj3+T
xeVWIkiF+WsLR8mBlDkmg8GUe5tajS5KuSREVv6dMFFlV45YYEbsFTJExtO2/CXi
Up7X0Lylizb7S7vY4sprWosy4Z/GcWoMePp3RHLsBDRl5uyMJbBoHtR6ITgj5E//
RHcMfnPWRUEfBT4dwF26alYkUaPX3U0Y2T4YMfuo+I6zmNthdS4usl46i3qJckek
tQWU0+/2cVbnTmd29W/KgNqjGd+eqpJCDe3oOtHFSdY80W2N8BQJfB0p3LIDo429
vI2LoLQgkwQ8OxIduRen1hfKFZoRlFX+S7fmYwLwCpeetzwvMUAj3vHGR1NZXA+4
3q3SajvxGmz69yaJLVG/d4YT+e+qU5Ll4kpfhLFXSiBgTvaC08U8zx9vggrxK9N5
f7sJHaTj2XIb9ZwdhzO4HNdZNM6Qp9ZFeDO1lVv8269cQBGNsQ27MzWnqe8sBZ7p
23iSx+w3klzpsMmzUt1LbAsMJa6esXaesZoFjYdl8OWkzC5v0H9s6JZwh83rd1oK
q98mH/zWfgXhESZDCpASW9hYvsjW3/GoH6YqL1YjBoYsfAclE1K4riYrZzMqfhWF
oGrC58DOFtfIlWeEnffaEe3GWkV1vRuOloYxDKHuAGa1R7jfZPyq3LupQ6OkrDn9
KUJufnheD1h0c3a6ZE7yr1Rhx1sPspepEj6Hz9JaY0eAoi8RMVIiAP6GFAGgIli/
Lep0bSBpETXligv9c0EbQ/WfR31/pXJuBlXc/zGBiADY1bn+Le95bpmkBxFRJI6e
EmPknW2hEdRDX/N++Q/MU+dGzhuQJ63+R6if2SrrlNVXOWbBCpft1vfhr2kYin5j
jJGakBJwt9QojoBSguhwMl6tZ3qyjEaZdj4fmV2X5BpvG2REOgq5RMxmAjA4q9xo
7m3VsyB6rfJngQ7zhC3vxvrLbeI/NssypD3z012PTOr5PDWg0E31qo3nyyJDHOhB
7upoQtugBYPplXfGrun2MLpBJwo/NLv3d4o1JedFVKEibavqTXj2DRd6n6FfzKxv
seaSoIhL769hDXedYIGczJbXkGnjs/jDBgtPwYqt+TkeElqAL0Iv/YwUdJ81RsHi
4D1+8/U4nE6etEOEUspM+YaV8dluWI7K0WbC6oblUvKbBlr2oX/iC8H5MGmPenB9
nqNligkWeUxjtpHuS7KawH/1EFNKHFPnQf6ET0JH00KaepzLuFgWATiXVKzeR2gO
yDvUUZNSr2xd//VV2IzuEmDvT1W+julRtHh0T085s45H4TQ4Hrg7+I3YNNq+98k0
mlF/j24f53kp8G1fleFtato+y/bUft6Z/UK/h/hXnQPQbS7CtTzQLLjuIlJQUB9Z
/AqcYf9DzbddXLHDqHqODZORTpo6+j+6HoPPwWmLG55Ieq1AbS2GrjL+mhmETSvD
T1Sf+JeTqsjMPYX9xQ0R8XWGSdb3J2RMtI42z154UMtW6WetgF0OMCiSuLlE440d
3v0RVl6gbDo5E1tY11fJohXZhiZCU4zIhRZp33mtp1FSzKyzdiR2DxhA5ip4QEcV
3tNzU6ywb7ps3TQ+nmz23ukRWhiXDQfu7HZMztNcywQhY+8f2SUnLe6RcMU7sVyv
JKYJcB1lZV610YxcKH8bAvITN2LCYitZDRnsbTBpSeyB/Hn8MIhyHGTIZumBBpVI
+tPe4gPVvQHqrm3OqDfEQVFA7kgbo74TXlDcx5P6Xtg1f2N71gvVGtUiNco4FoMJ
QuaUDb29omJzUsxRf8luT53cc+i+WI+iEUlHuug+OcMURhHnDWplYQUv7aIcSExt
1W/3fEqTk8I7LiZUihA7gwJiJmcde+acB7Oq0rXIal74jsMFUNuO755n6C6FU61D
5pKFZpbHraLAzDPuES1R+bctEEv+BMuQtOnHkFyrr1jFsvgklenaU3wEJdMoTn1z
VIwbperPCWqmv5HUARtGC7rrgrHSMI3Xi8PjCytFK3UOtz8EW3wiYcRTQYGlWOhN
8HbfQpzJG8CTiYWXCK5I1VsDWO9Ceqyibf3/+fJolxx/MAPEBeH1JKcYIVZI8Wk9
RAQkPic2XV4qEVmJXDQ40Xr81wfJtulooBoMuX//ZlQTmxWypJRl7jvPr8ZHFPx/
83mf5wuRGoqW64vxuXYG31w03npU+R7itMGVpBf87LL0rAK3C8ZaLNCNPdGY9M8j
2zAUA+6zYj/ZzBKkCXdfi8oTuKRMD44GNE3CFCtTbEIolBgLTtU3vf5uN1q665S7
Gz2n2LUc4m0bnNf127DsiUdiehB6hCuQz6eIyAYIKOBXWDXiOJ4/5e58DXQGoOtW
TIINx26Bpge40BeSiOTcy5WTaHYt9+QHnEjhw5zGS59vZvVYKU7TOYH57ace0sca
khDMs6IIk+cVoWbYe3wih56JVdjwcZjq/4I+FHzpIj4pgKDvsDHaRZdlP70T9lax
9E9VaQkCp2RoBDwqtYP0GoIW6sgHuvHV4IZcWw476Zql4V2qSHfM7xzlKYu9kIA7
POMzSMlP1QQ4poUrKXEindWeXUF+8/rCtz9LlVsPYkSbps8/V8V6ohFHcmrWwA4P
HzfNZR4KBWeA+TQ2VplMzqSpBSY8+0GpV5D5oHN0N3kCB1ohiUrhge9BPriZj8la
oc1x0F2QCqjO4Y5UtEWKPJBkXXbKJIgNhbNXtoIJtzXth31l8KqkGdypvGSJiZPo
cg+6idVKO5l0kvlY3AlYBlM4RjkcZn/YnB7YojOWIcxaZxX7/gntDvKFz7CI4J/c
jGbIWNWjVSTm4Y+NQT/QeRG3BcLAzKfuloAuG7Aa9Ohgu0M/h2s2+arZiX2Wb0Us
a/O7GLpyQ0bCuvtgDmjZMbzMUKGjU8C2o3ara3uZWQzvU3Mi/JXMMWE9p7xE/V42
dbI08YwNv5ApuElrvG0TMk4HpahYcCtkQBqHw/BbatF/Gv3NsCZBDPNA8jlwI/9r
YNdbTrhCQZKhMGy2m6puGj+cM2yTB3Kom9VZW73MPg+GkPscIwVZYr9PCZQik1Uu
md9F1xzwmdYEXiQNg3tmUDyV/RmaLBzw47nKB+KYPtM1GC91EK/iebNsairTMWOP
VSKv/YkEU0AgfxjGCFAgrgxr7Pan7Rv8+DOc84n/FTY5BdCOWKHFl8N5kxV5rUfk
em5CcUV+U37hCXJLLklyr+l//Upjh83y/tuntu3+kiPsdPU6nXY4rd+ZekgGkLHp
DyrZic1C3hXBfD4AddB0xkVEK0DcmJw0fmkeYbbEkRLW8Orr5b++R3YeW1GgmCoI
z+i6QsQpjhQWs9jQXB6Sn36bbuCIsJ4KgZJMZL0bkFtqKGBWnLM9Yn0agVCGYUYt
1YCrJlYzei7qRCrmJ7rFoMln+6tZwhthWl5Aoa8V85kDW8y9L+OwiOcIyKBsqLUn
xEszIbrI2S/ENSsiLMwsNUUbiKk35m6IZLgqFTNNJNXIjdBchCf79jQe3abgfJWv
4NyioLMUnYxwM0vYCqDlYEYJpMraz/gZgk8JqyhL+w6v1tCWgEytDhNlbSMXL6Ha
dCfWZnj7uPMmh6+UF3GxiyiZvECLtSEdq1hzg/fjlotu3MbmpzWphyeQdOc/lJc+
V0Sc/0y4BVio/q6vsnKj/ftRBiN9yJjSbdnkjyl0kzuefrN/vHo4Dus4KCMLSdJJ
4tvocG3ilUGjo717+PDs2eEwPxlM1tDzxKbAIsndWEwVGN84hBrMZz/L3zNLlOja
TRTlv/X0ykmFyA9D/Gs3vwv76GVbVlJcyLlqM/DL66XoygtQacNErwVz04hP46Y0
tQWYxNLgPC+uM4lLVFsa8YMiqx5YUPatvR1FAdXb9bcbqAtuXrGa7sEp4VUH4mhI
VbiVwC7qoLqWgLyXgTRWsW+R1/HARGmcB+rxnSWCDajr+ptBTxuj7qFeCWkbaY1s
rECrLoZwwQGy3jVAHCoQRN5Kd5qROzyUqW5exgXkM92UEztBHDsiL9VDCtg380Qz
jOBm+LxE9Rsx0Ls+4IWDD51/dDI/mgJ+9gzAU/lrUQ//NQ1oVr3aMs1WAXr5zNlk
kMMMUoP8NOGcSk1FOLzjfWHHywgghi3Mm+F0KbKw9v2mwR98yvc8f1Kjww9tlo+9
zc8HbGjLGti7pprxFnvvPdDiyLi92gr1Wwdg+GeM5knXJiAO/fcgGFCn9aECdBPr
suhdOxr4HL0PZoqjTYHFF9yGU/PG+yU+pLAaEUjQQjS/iyuz6agJSjw0nn8REOrP
iAlhm39C5qFDFNg9o9TnJB2JkKDHZ4JyGLzsdPwFpdxpgURUgWp8i8NqVBNaYD89
sHxpDzclZkvr2DugdPeSdtFcmSHiLrIxXNTB5GwwnPkS5kkBZAzPLPiKsA8ztkWg
8+cyu85QsouuDMeQGKAW1kXH8U1rmCYG0jG6rGYStABEtZr9Zg+nHiB9LD3qIJnG
SeOHq9HUyzMRKbKdmUv6stgEdD5qPLaACbzt3z4v/LQLGyxkj9VNxTYB/kczwmBr
M0FtbfhC/77gC85wnJQJF3dyXOnN4EWPezmcyZdXIR3/gr4CJvv6kvDGd/BjbIxY
VGQ5BKS0ZwDZzNisV6ncMXEgXoBBzIBUdcyBgjdOOME+2/yVZlozab8sx1TW96pd
vzQ9sqBsMf10eheotu9+9SmiHgWniZKf7+7rzhJzfrFfVdwHmd2BYRxKv89jTbcM
l28HtlUe8HLKxx2X2lPtDKVco0xIaHf1bPfwOhQ+RPc=
`pragma protect end_protected
