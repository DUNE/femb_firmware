// Copyright (C) 1991-2014 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1.4
// ALTERA_TIMESTAMP:Thu Mar 13 15:23:41 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
K+VREjMSYN5SWJPZsdlBTnx7u2tVIjZaIwE1lSXwcuX7diRRiK0gju3Md17AKp/j
fENOXEsyQjZs9ZgdUSQuClld4qGKubCB5anKAsmMJzawTsIcWn1F6l+2ydCSq10m
PPD5IZbvH8YTveHOMDXi8lgiRz59nCXL1+l/BgcOKxg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5488)
G1OYnaop3v0NipYtFy7v0hqLCiECWegdzsUMaQ9Wi8q9Y7NSW7dHMaS6XNz5XHuP
CLE5LUQBGtfLfUqEGZBNtNN9Zbt1n3LxgBhdXELxovn7DnEFbyK/OqakqjFrjxfv
TG97bwNIhudZYMtavYvH5WjPYWEczO5/eC94VQ8DBEg3B1OGaNGQD4E9CxHflNPW
62NUYZOAwkPHq5veY/qBPtsHJiesY2HIAfFXbkF2xToCWtX2mDC38lO1Nc2M1RwU
5qQaEcAOXLfBPSSZIUJVcumMLGB3bCuOm+FS6vx8uSE+KVyBj0tzadELSahbheLP
x1ZQ67K7PES4y9Xe2nlrp1bLIpEmsTSxu9MCV0pULsetsUErUJ8YSm95lnmhZ36h
kExbdbD+iHiQJbmGQQ/DCJdU/bs3ALb+YtufF0RqEZboPg47UMu+eCcYH8wejKP4
Wdx4+7d0m9osuR0TL07QYwx01t6CFSgALZlBWA3jg3T1R10fWJpcOG2/B/XrVr3l
t8JM6P5IoJdd1OYXvMboTc3hEiSNEwv7VbSg0tNj0as8xFKTFH0U20fLzrnbL6+g
fsEHXa8QFmEfzPWZK5RxfQudTbydkYzbcqtb5Y/XR6ksMHl2w5TCUaD2z97l9NaO
SlRkPuuKaNrEG9LdOELuICwtTutRNcj3ap9Z58R+cVcqOS+YWCOWGaM5ZinJbaa7
cVlp3Upwxvl23Cs6AEvtpTqqdcIb43ynuQjuthM19Ailb4YwJbHM67ojrGpy4liw
tHn8ncqPhLPwKs8eY1Hw6Oh97PooFKuI6sRogDuimmQ0be5Dj+VZe5YEUFvVkC63
Y2XV82DgjTvHpjReBUPI+407+LmtuPvTRNoQNWzanef/2+7sQYOB9z4U09jqCZ+g
jJemJnzcHq/1nbYSm6eV2P4sTUv1KXv1iT6pTs4ozjjQ+Y9OYZBpSSTJ4qZoy0IM
zzNxdPiM4o+oVkz8aptbyS7TIpvXu7hjUlAiDpTSwAXelw89oFGls8f9sEs7xAEf
GeHxld/a6x3I+JvfDOTCo5L4GdPRA3ChZMvHs1wUr/h+O7njQhjqp6NK7IzTv0lh
ODF1mmi1K2oKT1kJTdC9I7WZrFgBvPzT6mCMRUZgrp5Kt4MwtNlcRw9X3Bh3koHP
3E2mTmtj4ZZu2OkFbueARpB3xQrcPr0jdMca9L+6o6NTx2mXELwUhrGMkQS/WMm8
KRLGe1ivg/JWvfelEb9MppkZ1/zak+/KINnecnry2cHoUJcdvGhJno6Hiq8OdVKN
04bSZ36I77ayPGSKev+sPQzEbzDMD6sO3JBhfB/V9Sdf1tIPkb56cHAdVkysgBel
30ZnUyWhTTum+nI3n2ydnyZr+y/R9q1dTwMSZfwDEkU23GQMaphnVRHhG5mpXifc
artHBSgjxVzKT2UaHDalxkluJoimV1WbOa4Iuly2RfY5xfApdKo+0lk7d7i88pxP
NTBSTK4njmIT8fAuUVTNPAQsFvMEno7Wyw1TD3WRAnnsGxrhuIzd93FRTMlZkKIt
CwpCz2OQVrQp+qxiDKr+TnYVIaqtrF+G2Bg/MnlNm+aKCBPZDDMWqPIBLr+LIRAI
TDznfIa0UazVgx4ovpVTej2E2HB75d6NfPLsfPXtwDK35m2MyDBa5GDY8nz1XCGo
4iJyxfj/TWXGoTXKqOCDc+ugJMXhJhp59/nbBXimixT2uC9iNtLIQkjToeW75AMU
4hIlhceiPmN5AG7X9ENd4CjDrOvWXyFxb8s1KlIdPkQh36FteYEA2VB3y/9wm385
gQgUS7df2Dd3zQiyKcli6WVfK/fovmjIXtfjWlQQjECaAfmuQOKTLxFYL1c8Ev9z
UtvouE2nbSXp+cNVsGRE0IEyKLvoGtAzw+GJrhLxyANsNLImE58s6SyH/97S736m
y6PbJwCidqswba4PwwJpbMcfN/SbuFJGNSvxEfX/vEhHt9WK7K0BDX6ZdlfatXLu
htGZENILvsxyYpg2kuSTPa758tRk7DMfB++qU3AUzU1QNir6HInbWHVjaSBlxsgP
ApKKdsai3BWcCa2qZ8b84UL4lAPj78vLQ2QPwOiL2d828LmTqALW8vu12N8bOFga
1p8FsDXfTPQISmATGFmtTZw5cb37dgHqznyadpXTiqH0xWvua1WYuTN2r2Q5OiWs
pAhwlVbjkleyEeBoR+9dU3/gJd4iAcFAeJwvkgeIMmqbyqXkyKmmNSotLgHcz38I
NL761RdWU3lCdM8jVU24+39H3Ugg9vBe8ZijUeKkrtXzTY52F8yPotrm2lK/KXYa
JoV/J/nVnbyvJcGGw8jxiC3oK+gQiMbjttqePb3x1kv8Vcku67/Xr73OZFwOtfq9
HkkIPlSLQrBdFoVL0M6ZNWYFDBoEJqVsw4UT6PC8ssa3vhBKqHZXA+BtmmpCsO9D
PG6mUUVTjfLxjy5O+wKDz53ywMB4XcQ3uvRzGMp2QigZOHo7OtCRkY5jXeQ+1s3M
8GcLjNokTFWDEwXng41+MAf2FmwZUolY8BviUvFV4WJqueOKsEQvsZou+9kikeKh
u0l9gk/dPhdA1MIqIvcOs9Ghn8MkmwZRypZ2uuLOJBS97RuSjUQTVWRgobJzYQSr
Bf6N8UT9FH0wEuKBIa24VnmuEcaDuQQrD1z5zF8lKQCnMlkhtIdyohx5f+v6cVVs
2U/eJCymR2V0m/6nl2kWA/pKFh59JB/K4qQRkaBmARot3zJl5FhhwqRLrhORjogJ
WEWE+c3LOjche3P68gAa70d5Pj3QcmURQfsSDDY5xdm20+09ovMZ1aQ042ETaJOT
G+qzfw+ptaUI4UdKhcwRVXQzhR20ajwwCnvWE2PT7B+UBzF5txduDcSglB5sIFq1
RWBDfHi60G9T+VPf6RRHr/yxdIWWJK6URIhUPzci5uVGwh3ftEHGqHUj0En5YOxM
lwHmAn6Vc0aKfCwP2IMv7TfQo1idJqR/mEJ5T18zYWc1WG7abOEjWUKG8laMCn2v
YpxK18/+Xkak/k17zudtu+/w/b0q5ElPAjaCRIg/ANiXlkCFHAn8sVOx1fdLW7Ru
T66PMe3KwxLF7h1OkFwQtFozJDv3d0ZQeUd0P617CxjK53DRXAeqpoJDPhtzVeHN
ncVnGKwMhcy9JmVksC7xkb7W7jNjfLShUsuMLQj5VzDQbwnSwAlkGul9xGJvJtNg
s9EpRP4BK2Z3USz9tqU0SdoYQiTXTqHLArBhGkIuz9WhiGTpEIKuKnUutJJDMZIU
a0LRmKrXfsCHuLrmdNL69hLNzTM/3FrOk5DP3/dhpjUYV57d5SFbPKbsERfraI4v
NsETXK57iTEm6dfkr5U/pRh24PbAdr169DafJQSJzcoumM4Jl1wcfH85rikpAW6u
tbSE6X6ZHJ+71uMrzTJ/Z3Dmefx7Bq8HMWWPxPOePIzlY9fdpu9RvwlEoYxybp29
8o94qaFPkkNx7m8w2k3jEr2FSE3liPrCoYdIPCIqXaYopk30hEoKCXz7lDNLoEdK
8aDmrdSE0etjN/QbGvIilRzGrJbS+roxFQvUaVnp0JO6omRC+IfL6W91CSGqziIH
lIhB2AmoyqmSNtrKuLRABkENO6aUYUTIooJDj5SXi7aQZ6+YtG7g4XNbVH1JNQgZ
7glaf0rufXhH+/Zd6cQB6RjkJgdkrcqMxAiFUTUQ8Fe9gu6ZKPkG0ryqdzpXYNCh
/rSsn16SBCLu3HVii30pKxeXUt4SQMPIORjDJAOjzrJkGyxtiZNA7HO6fByRZO+V
ztSKj6okmtC5bxAop0qSiFdXwdWSlB/vV9CNcJyZHl+eKTe/meLINhEfLeqXl409
m7jUFhGCX/uNpe1iaZ/X7tAnq9B4tNjQEEe+k4DNSdcgP95QWh4l/B0ugBbayKI2
MPgeELlqtWCEtQyicrMQOqt1kpOELpiqZEh4dJmVATgXsk/OfSHWrM3AqGlFhaRn
G2dgI4k2Igqa1XdoGGIHdkvIUkTsZ8tLKFsFimKNcdF1nvPVz98cdPKDx9NHLORr
HTxVt3mJd1qZcQuZhJhT+PBXPmdgd7f0zE4grvrRTsF9Z9eYEjkARLGJL99YXSIO
mG4XEk+SHBpwy76SYzf1rYi+t+8NNsjPjqcf7b4ZCMUldEn1S3eBFKRZSqFH9e7H
s1duO9B1SQu11O7HIx4cJKrhyIWZGL0H+tJCoIXvOSztb3Srh1vdYWvfiZ7/LLzB
v7pX0JgU7wvy2GMpPneER0ssCTeoJNyF1dwYTdwZTmQaocUswK/d4bJYWWXkn6eM
gSWaroRstwoR9h941wGJJ35iijF6foWxJxJRwrQnpoGgtoVTze/f28x0ONUC6EPV
M+VMwvVCPa1R+T+4wLG8K7GBbGv7RvnTRawkDZ3PJjLYs1BvngHWIYcavb2EdMI3
4jcYD4qpM16hMYYIBQ851Uvvs2Wu5QNYiZbd1W3dgwgDO1LBWjARgFDvHecirotc
rLSrNxUoEW+eEkjAfJMjHRkVgKV54OKL2/98AWIyqdghqmHcATkwPuQJBPqvHYCA
jN2w2tAvgear8FAGTT/fRW6d4YdOIg7Ft5ECd2rI1v5d6y35tWMYSJMSuvOqM0Cv
wWo7HWp7Vj4incvA8SR3NrRptGCp1qz10Z0FAclTnJXGZ4ZrZgxvjuGDdd6IGhqp
zZgBl3od1Uc8RV+w3CnS0bMoFBg3C4MLptHzg+helw0rm1K7ofPXwq4c5F/DqAU5
7d3ev/+pw2fVU0bWiHaq+ynKdx28Iwcoy6j4UfYh9tRe+g+xcD2P1EFws/nCO+0D
ThXroPUD4sqJLrY0VthWyYKIL+90DYm+uiaqv2WAFmTKfIGzeM7i9+sqTKsqpqU3
NVL2kXuILpv4zBaWOQqEDQLISnipY/oGi+I5nhpMrNvlAXJmVfxJXM8KAw+41i7I
MvPZoJwrNtGUOAsJXdu6GCNYySqdY4DSGqSH/EtvD1GUJ8/wyi3YqIPDt6Ge0bjj
tOZq8uyB9j9OeT+OOHJYri0vqs9dNTPMRlGh28ERw13DvF/vPK4Wcyw5e5v/yQPh
TesYBebraz7AAvD4UPIl1gNluPa/aux+So7xNi7YrupyP3+BuDYjJqj4TP4IGhfq
AhbbkMYRfuNW5cr3DbibYVhbbMjCk19tXP7CZUY1ObqlvJKMJKyK5NKFPa03FOQv
2UdaGA4NDDTfEEaU8uMQzuer+oq9XZlBEGUAgl3yusOAyssuAQv9iiMQedSOcgXR
IzwNR4Vczr7Cp2nfHOoKuVAU6XtaGeBxkEiYMGdXyBAM69tXfbMoTYitYyTQRQyu
TguYN0S6U/qx+l0krOQ5rJFkscoryiLOqCOFkaRf3TLPJCeRrn44zq9PcmLD9Tpb
qthYtNTBxpaYOil8474CDfkx8jlnl2Tp6uEfVg5t6cwketVEjPopxP8MoRmC/J06
y56076mGiUNIOgvLsTlq1MEcBcpxyT0Idy262sdcMltcdqkPQoFdbFyq2CTJLjA+
sLJJcoiJg3dg32ctvP2Zs51EGhanbGhh/nNZMLbAeGs/o2G8bNL7lRC8UvWgnY6X
0XIBFgia3CCVCNWe+hwQG0yH2mniWuMY90ON31a1D9kAtV8533chswQG9aKLjTTb
EiUflPMvBZCbe0dkEL/9TWaTt2aDuaIFekL79REu3rH4KrGYBMCmOeojUrsOZUno
//y+G0WtGRtCkZksDQvzdQjumzK905kNPG+mKyR+WkrVvHAf8V2fb/oh3DEkR5uB
3FbcpmOfh6iwdlpu5y5poMHXzZzyD/3pXiOkIa4a+A58RxrUZx0ajYBclMovpyXX
+cDAHG7/m0Txv1c2mO6+vJvca2CAdNKpf6yHS1uTiQCe02eQAPePhEqdM/Fd18mc
b6qcBpuISiITM7GBkHTR5+PFs5P2Rj94KP4C8uGbmenlCDhmRXhXPZlWT29DCU6+
1jNYzAdRRstgxx/o4qYJqJqu+CAeMG3YYgEF1enjXxiVbRWwNJOmzeozrFHwltRG
/PhFEzwRLVd6vGO/YtMmP8GvIqHCW+kp7a4bX+ibVX/OblDWedY3QafHeHPaWSFt
rzSPedxQLKyxfvo43u0TWob/p6wFoF8pzzFtD5n+rxek9DCJE1Uldq1vItdUhw6T
vUJHrca5MrSqpME0KKB1hC7eL4LcYBJeWLmOn7QeHhhSMbaMIXKS3kzRw/R8+9XO
3QKqn/lI/NlRtlx9v+VlUc1SCsj2tJFfbhs8AJJh2B/A2ucXGcioLkgVA12z4BmQ
TuevDCTCFJ/O1Cwcs2l45feG1pnTu5xkMQLA7oxRnh3IMO487ThEx7CbKKr7N75f
UO8Ut+2P1eGZYJ6kf3edtBBuhjLpE2+Fjcr3kwYbAeshCy6KQGGHsLpCsMlyQ581
Jg0kKP6ZG1NGUQ3KdhV7rWIE3GugQTZhPtARXuzOob8uh6YsCgAWPnKx51aJ0ORt
qkWjC2ZuBzuh/9qpv+23FiKyRng74gOpNG1L83IvdffNWyf4CZQ4KsLYRdNcwewg
M+XZOqThxiwpA9oIBxW6V5vI8OyodfXR3VFrrlW+Aj6pl5oiQcG7LPS3WLrzKXNW
PrbQEEC+4oWIy3C+mAnK0TruTWZAi4VomwBTP4KuZHwoSUuLdJqizGK/t/li0gec
AvBJrxycqrJGyjUTIQFIzgtdUevuIFTm1Pe//Hyf+/Q/jaY+Y5Fa+xiNgMPzel1h
vsMKq4iMherQHYJTIvSuA/fa3iw0uVGkBmt2d32yJQ5FHRz02SZC4zjJI3dsdw4x
Y5DpeSveERuffL+r2B7GYxwwFyexHKITJZjenTeJYKPWK+dM2UO6pyRMIkSbTt9T
00WdcsVzMBCzjiUMKDBXd28fpqSTaRBh5zRgGhKBkVF6kXn65sxST9oAjwAjfBnw
MoGQgMJzE1B16/I5qM8D8dMp1IVsg50YZ5APkUIcDTSDAiAkAui0Pf++mCJsY3m0
SW0P8m1OHntkbFXzjGB2fQ+JLkO5/obXVRgU39v7oxs0gb6XUhTZZgLUiAeYx5Vz
5LpxQZNQsTCICmrMFvm58DpiTzWdt6w9mLCMl1QFvPWj/rDci//u9qRmSh8xdbH0
yAY8q+avIHnqiDWkWaDox+9FSU0ow9/hA/SEyse87hy8rTrq1OpbzHBH5bq7TIPH
wU86uRRMrhc70bMMu0iQiQq4zD3uCKGGGvg4L22UnNBv9ay59o8dmxyg8u2VpRxl
B5/To00LwEXOoAqrh9jNy5PpJIpEJkhvARBcGlll+qmzWPnXZO8O6ATl8Ad4X5pW
7BCCPBfDpBm4+g+poAq1bg==
`pragma protect end_protected
