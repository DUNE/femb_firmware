-- megafunction wizard: %ALTGX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: alt_c3gxb 

-- ============================================================
-- File Name: ALTGX_TX.vhd
-- Megafunction Name(s):
-- 			alt_c3gxb
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 16.1.0 Build 196 10/24/2016 SJ Standard Edition
-- ************************************************************


--Copyright (C) 2016  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Intel and sold by Intel or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


--alt_c3gxb CBX_AUTO_BLACKBOX="ALL" device_family="Cyclone IV GX" effective_data_rate="1280 Mbps" gxb_powerdown_width=1 loopback_mode="none" number_of_channels=4 number_of_quads=1 operation_mode="tx" pll_bandwidth_type="auto" pll_control_width=1 pll_divide_by="5" pll_inclk_period=10000 pll_multiply_by="32" pll_pfd_fb_mode="internal" preemphasis_ctrl_1stposttap_setting=0 protocol="basic" reconfig_dprio_mode=0 rx_enable_second_order_loop="false" rx_loop_1_digital_filter=8 transmitter_termination="OCT_100_OHMS" tx_8b_10b_mode="normal" tx_allow_polarity_inversion="false" tx_bitslip_enable="false" tx_channel_width=16 tx_clkout_width=4 tx_common_mode="0.65v" tx_datapath_low_latency_mode="false" tx_digitalreset_port_width=4 tx_dwidth_factor=2 tx_enable_bit_reversal="false" tx_enable_self_test_mode="false" tx_flip_tx_in="false" tx_force_disparity_mode="false" tx_slew_rate="low" tx_transmit_protocol="basic" tx_use_coreclk="false" tx_use_double_data_mode="true" tx_use_external_termination="false" use_calibration_block="true" vod_ctrl_setting=6 cal_blk_clk pll_areset pll_inclk pll_locked tx_clkout tx_ctrlenable tx_datain tx_dataout tx_digitalreset intended_device_family="Cyclone IV GX"
--VERSION_BEGIN 16.1 cbx_alt_c3gxb 2016:10:24:15:04:16:SJ cbx_altclkbuf 2016:10:24:15:04:16:SJ cbx_altiobuf_bidir 2016:10:24:15:04:16:SJ cbx_altiobuf_in 2016:10:24:15:04:16:SJ cbx_altiobuf_out 2016:10:24:15:04:16:SJ cbx_altpll 2016:10:24:15:04:16:SJ cbx_cycloneii 2016:10:24:15:04:16:SJ cbx_lpm_add_sub 2016:10:24:15:04:16:SJ cbx_lpm_compare 2016:10:24:15:04:16:SJ cbx_lpm_counter 2016:10:24:15:04:16:SJ cbx_lpm_decode 2016:10:24:15:04:16:SJ cbx_lpm_mux 2016:10:24:15:04:16:SJ cbx_mgl 2016:10:24:15:05:03:SJ cbx_nadder 2016:10:24:15:04:16:SJ cbx_stingray 2016:10:24:15:04:16:SJ cbx_stratix 2016:10:24:15:04:16:SJ cbx_stratixii 2016:10:24:15:04:16:SJ cbx_stratixiii 2016:10:24:15:04:16:SJ cbx_stratixv 2016:10:24:15:04:16:SJ cbx_util_mgl 2016:10:24:15:04:16:SJ  VERSION_END

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY cycloneiv_hssi;
 USE cycloneiv_hssi.all;

--synthesis_resources = altpll 1 cycloneiv_hssi_calibration_block 1 cycloneiv_hssi_cmu 1 cycloneiv_hssi_tx_pcs 4 cycloneiv_hssi_tx_pma 4 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ALTGX_TX_alt_c3gxb IS 
	 GENERIC 
	 (
		starting_channel_number	:	NATURAL := 0
	 );
	 PORT 
	 ( 
		 cal_blk_clk	:	IN  STD_LOGIC := '0';
		 pll_areset	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '0');
		 pll_inclk	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 pll_locked	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 tx_clkout	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 tx_ctrlenable	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 tx_datain	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0) := (OTHERS => '0');
		 tx_dataout	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 tx_digitalreset	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0');
		 tx_seriallpbkout	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END ALTGX_TX_alt_c3gxb;

 ARCHITECTURE RTL OF ALTGX_TX_alt_c3gxb IS

	 SIGNAL  wire_pll0_areset	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_pll_areset_range39w40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pll0_clk	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_pll0_fref	:	STD_LOGIC;
	 SIGNAL  wire_pll0_icdrclk	:	STD_LOGIC;
	 SIGNAL  wire_pll0_inclk	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_pll0_locked	:	STD_LOGIC;
	 SIGNAL  wire_cal_blk0_nonusertocmu	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_adet	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_quadresetout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_rdalign	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxctrl	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxdatain	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxdatavalid	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxrunningdisp	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_syncstatus	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txanalogresetout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txctrl	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdatain	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdetectrxpowerdown	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdigitalreset	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdigitalresetout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdividerpowerdown	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txobpowerdown	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_clkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs0_ctrlenable	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_datain	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_datainfull	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_dataout	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_forcedisp	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_powerdn	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_revparallelfdbk	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_txdetectrx	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs1_clkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs1_ctrlenable	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs1_datain	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs1_datainfull	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs1_dataout	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs1_forcedisp	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs1_powerdn	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs1_revparallelfdbk	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs1_txdetectrx	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs2_clkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs2_ctrlenable	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs2_datain	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs2_datainfull	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs2_dataout	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs2_forcedisp	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs2_powerdn	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs2_revparallelfdbk	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs2_txdetectrx	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs3_clkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs3_ctrlenable	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs3_datain	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs3_datainfull	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs3_dataout	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs3_forcedisp	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs3_powerdn	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs3_revparallelfdbk	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs3_txdetectrx	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma0_clockout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma0_datain	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_dataout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma0_seriallpbkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma1_clockout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma1_datain	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pma1_dataout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma1_seriallpbkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma2_clockout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma2_datain	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pma2_dataout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma2_seriallpbkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma3_clockout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma3_datain	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pma3_dataout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma3_seriallpbkout	:	STD_LOGIC;
	 SIGNAL  cal_blk_powerdown	:	STD_LOGIC;
	 SIGNAL  cent_unit_quadresetout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  cent_unit_txdetectrxpowerdn :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  cent_unit_txdividerpowerdown :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  cent_unit_txobpowerdn :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  gxb_powerdown	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  nonusertocmu_out :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  pll_powerdown	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  reconfig_clk	:	STD_LOGIC;
	 SIGNAL  tx_analogreset_out :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_clkout_int_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_core_clkout_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_coreclk_in :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_datain_wire :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  tx_dataout_pcs_to_pma :	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  tx_diagnosticlpbkin :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_digitalreset_in :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_digitalreset_out :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_forcedisp_wire :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  tx_invpolarity	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_localrefclk :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_phfiforeset	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_pma_fastrefclk0in :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_pma_refclk0in :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_pma_refclk0inpulse :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  txdataout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  txdetectrxout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 COMPONENT  altpll
	 GENERIC 
	 (
		bandwidth_type	:	STRING := "AUTO";
		clk0_divide_by	:	NATURAL := 1;
		clk0_multiply_by	:	NATURAL := 1;
		clk1_divide_by	:	NATURAL := 1;
		clk1_multiply_by	:	NATURAL := 1;
		clk2_divide_by	:	NATURAL := 1;
		clk2_duty_cycle	:	NATURAL := 50;
		clk2_multiply_by	:	NATURAL := 1;
		DPA_DIVIDE_BY	:	NATURAL := 1;
		DPA_MULTIPLY_BY	:	NATURAL := 0;
		inclk0_input_frequency	:	NATURAL := 0;
		operation_mode	:	STRING := "normal";
		INTENDED_DEVICE_FAMILY	:	STRING := "Cyclone IV GX"
	 );
	 PORT
	 ( 
		areset	:	IN  STD_LOGIC := '0';
		clk	:	OUT  STD_LOGIC_VECTOR(5 DOWNTO 0);
		fref	:	OUT  STD_LOGIC;
		icdrclk	:	OUT  STD_LOGIC;
		inclk	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		locked	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  cycloneiv_hssi_calibration_block
	 GENERIC 
	 (
		cont_cal_mode	:	STRING := "false";
		enable_rx_cal_tw	:	STRING := "false";
		enable_tx_cal_tw	:	STRING := "false";
		rtest	:	STRING := "false";
		rx_cal_wt_value	:	NATURAL := 0;
		send_rx_cal_status	:	STRING := "false";
		tx_cal_wt_value	:	NATURAL := 1;
		lpm_type	:	STRING := "cycloneiv_hssi_calibration_block"
	 );
	 PORT
	 ( 
		calibrationstatus	:	OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		clk	:	IN STD_LOGIC := '0';
		nonusertocmu	:	OUT STD_LOGIC;
		powerdn	:	IN STD_LOGIC := '0';
		testctrl	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  cycloneiv_hssi_cmu
	 GENERIC 
	 (
		auto_spd_deassert_ph_fifo_rst_count	:	NATURAL := 0;
		auto_spd_phystatus_notify_count	:	NATURAL := 0;
		coreclk_out_gated_by_quad_reset	:	STRING := "false";
		devaddr	:	NATURAL := 1;
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		in_xaui_mode	:	STRING := "false";
		portaddr	:	NATURAL := 1;
		rx0_channel_bonding	:	STRING := "none";
		rx0_clk1_mux_select	:	STRING := "recovered clock";
		rx0_clk2_mux_select	:	STRING := "recovered clock";
		rx0_clk_pd_enable	:	STRING := "false";
		rx0_logical_to_physical_mapping	:	NATURAL := 0;
		rx0_ph_fifo_reg_mode	:	STRING := "false";
		rx0_ph_fifo_reset_enable	:	STRING := "false";
		rx0_ph_fifo_user_ctrl_enable	:	STRING := "false";
		rx0_rd_clk_mux_select	:	STRING := "int clock";
		rx0_recovered_clk_mux_select	:	STRING := "recovered clock";
		rx0_reset_clock_output_during_digital_reset	:	STRING := "false";
		rx0_use_double_data_mode	:	STRING := "false";
		rx1_logical_to_physical_mapping	:	NATURAL := 1;
		rx2_logical_to_physical_mapping	:	NATURAL := 2;
		rx3_logical_to_physical_mapping	:	NATURAL := 3;
		rx_xaui_sm_backward_compatible_enable	:	STRING := "false";
		select_refclk_dig	:	STRING := "false";
		tx0_channel_bonding	:	STRING := "none";
		tx0_clk_pd_enable	:	STRING := "false";
		tx0_logical_to_physical_mapping	:	NATURAL := 0;
		tx0_ph_fifo_reset_enable	:	STRING := "false";
		tx0_ph_fifo_user_ctrl_enable	:	STRING := "false";
		tx0_rd_clk_mux_select	:	STRING := "local";
		tx0_reset_clock_output_during_digital_reset	:	STRING := "false";
		tx0_use_double_data_mode	:	STRING := "false";
		tx0_wr_clk_mux_select	:	STRING := "int_clk";
		tx1_logical_to_physical_mapping	:	NATURAL := 1;
		tx2_logical_to_physical_mapping	:	NATURAL := 2;
		tx3_logical_to_physical_mapping	:	NATURAL := 3;
		tx_xaui_sm_backward_compatible_enable	:	STRING := "false";
		use_coreclk_out_post_divider	:	STRING := "false";
		use_deskew_fifo	:	STRING := "false";
		lpm_type	:	STRING := "cycloneiv_hssi_cmu"
	 );
	 PORT
	 ( 
		adet	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		alignstatus	:	OUT STD_LOGIC;
		coreclkout	:	OUT STD_LOGIC;
		digitaltestout	:	OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		dpclk	:	IN STD_LOGIC := '0';
		dpriodisable	:	IN STD_LOGIC := '1';
		dpriodisableout	:	OUT STD_LOGIC;
		dprioin	:	IN STD_LOGIC := '0';
		dprioload	:	IN STD_LOGIC := '0';
		dpriooe	:	OUT STD_LOGIC;
		dprioout	:	OUT STD_LOGIC;
		enabledeskew	:	OUT STD_LOGIC;
		fiforesetrd	:	OUT STD_LOGIC;
		fixedclk	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		nonuserfromcal	:	IN STD_LOGIC := '0';
		pmacramtest	:	IN STD_LOGIC := '0';
		quadreset	:	IN STD_LOGIC := '0';
		quadresetout	:	OUT STD_LOGIC;
		rdalign	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rdenablesync	:	IN STD_LOGIC := '1';
		recovclk	:	IN STD_LOGIC := '0';
		refclkdig	:	IN STD_LOGIC := '0';
		refclkout	:	OUT STD_LOGIC;
		rxanalogreset	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rxanalogresetout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxcoreclk	:	IN STD_LOGIC := '0';
		rxcrupowerdown	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxctrl	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rxctrlout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxdatain	:	IN STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
		rxdataout	:	OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		rxdatavalid	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rxdigitalreset	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rxdigitalresetout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxibpowerdown	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxpcsdprioin	:	IN STD_LOGIC_VECTOR(1599 DOWNTO 0) := (OTHERS => '0');
		rxpcsdprioout	:	OUT STD_LOGIC_VECTOR(1599 DOWNTO 0);
		rxphfifordenable	:	IN STD_LOGIC := '1';
		rxphfiforeset	:	IN STD_LOGIC := '0';
		rxphfifowrdisable	:	IN STD_LOGIC := '0';
		rxphfifox4byteselout	:	OUT STD_LOGIC;
		rxphfifox4rdenableout	:	OUT STD_LOGIC;
		rxphfifox4wrclkout	:	OUT STD_LOGIC;
		rxphfifox4wrenableout	:	OUT STD_LOGIC;
		rxpmadprioin	:	IN STD_LOGIC_VECTOR(1199 DOWNTO 0) := (OTHERS => '0');
		rxpmadprioout	:	OUT STD_LOGIC_VECTOR(1199 DOWNTO 0);
		rxpowerdown	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rxrunningdisp	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		scanclk	:	IN STD_LOGIC := '0';
		scanmode	:	IN STD_LOGIC := '0';
		scanshift	:	IN STD_LOGIC := '0';
		syncstatus	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		testin	:	IN STD_LOGIC_VECTOR(1999 DOWNTO 0) := (OTHERS => '0');
		testout	:	OUT STD_LOGIC_VECTOR(2399 DOWNTO 0);
		txanalogresetout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		txclk	:	IN STD_LOGIC := '0';
		txcoreclk	:	IN STD_LOGIC := '0';
		txctrl	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		txctrlout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		txdatain	:	IN STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
		txdataout	:	OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		txdetectrxpowerdown	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		txdigitalreset	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		txdigitalresetout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		txdividerpowerdown	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		txobpowerdown	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		txpcsdprioin	:	IN STD_LOGIC_VECTOR(599 DOWNTO 0) := (OTHERS => '0');
		txpcsdprioout	:	OUT STD_LOGIC_VECTOR(599 DOWNTO 0);
		txphfiforddisable	:	IN STD_LOGIC := '0';
		txphfiforeset	:	IN STD_LOGIC := '0';
		txphfifowrenable	:	IN STD_LOGIC := '0';
		txphfifox4byteselout	:	OUT STD_LOGIC;
		txphfifox4rdclkout	:	OUT STD_LOGIC;
		txphfifox4rdenableout	:	OUT STD_LOGIC;
		txphfifox4wrenableout	:	OUT STD_LOGIC;
		txpmadprioin	:	IN STD_LOGIC_VECTOR(1199 DOWNTO 0) := (OTHERS => '0');
		txpmadprioout	:	OUT STD_LOGIC_VECTOR(1199 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  cycloneiv_hssi_tx_pcs
	 GENERIC 
	 (
		allow_polarity_inversion	:	STRING := "false";
		bitslip_enable	:	STRING := "false";
		channel_bonding	:	STRING := "none";
		channel_number	:	NATURAL := 0;
		channel_width	:	NATURAL := 8;
		core_clock_0ppm	:	STRING := "false";
		datapath_low_latency_mode	:	STRING := "false";
		datapath_protocol	:	STRING := "basic";
		disable_ph_low_latency_mode	:	STRING := "false";
		disparity_mode	:	STRING := "none";
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		elec_idle_delay	:	NATURAL := 3;
		enable_bit_reversal	:	STRING := "false";
		enable_idle_selection	:	STRING := "false";
		enable_phfifo_bypass	:	STRING := "false";
		enable_reverse_parallel_loopback	:	STRING := "false";
		enable_self_test_mode	:	STRING := "false";
		enc_8b_10b_compatibility_mode	:	STRING := "false";
		enc_8b_10b_mode	:	STRING := "none";
		force_echar	:	STRING := "false";
		force_kchar	:	STRING := "false";
		hip_enable	:	STRING := "false";
		logical_channel_address	:	NATURAL := 0;
		ph_fifo_reg_mode	:	STRING := "false";
		ph_fifo_reset_enable	:	STRING := "false";
		ph_fifo_user_ctrl_enable	:	STRING := "false";
		pipe_voltage_swing_control	:	STRING := "false";
		prbs_cid_pattern	:	STRING := "false";
		prbs_cid_pattern_length	:	NATURAL := 0;
		protocol_hint	:	STRING := "basic";
		refclk_select	:	STRING := "local";
		reset_clock_output_during_digital_reset	:	STRING := "false";
		self_test_mode	:	STRING := "crpat";
		use_double_data_mode	:	STRING := "false";
		wr_clk_mux_select	:	STRING := "int_clk";
		lpm_type	:	STRING := "cycloneiv_hssi_tx_pcs"
	 );
	 PORT
	 ( 
		bitslipboundaryselect	:	IN STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
		clkout	:	OUT STD_LOGIC;
		coreclk	:	IN STD_LOGIC := '0';
		coreclkout	:	OUT STD_LOGIC;
		ctrlenable	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		datain	:	IN STD_LOGIC_VECTOR(19 DOWNTO 0) := (OTHERS => '0');
		datainfull	:	IN STD_LOGIC_VECTOR(21 DOWNTO 0) := (OTHERS => '0');
		dataout	:	OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		detectrxloop	:	IN STD_LOGIC := '0';
		digitalreset	:	IN STD_LOGIC := '0';
		dispval	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		dpriodisable	:	IN STD_LOGIC := '1';
		dprioin	:	IN STD_LOGIC_VECTOR(149 DOWNTO 0) := (OTHERS => '0');
		dprioout	:	OUT STD_LOGIC_VECTOR(149 DOWNTO 0);
		elecidleinfersel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		enrevparallellpbk	:	IN STD_LOGIC := '0';
		forcedisp	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		forceelecidle	:	IN STD_LOGIC := '0';
		forceelecidleout	:	OUT STD_LOGIC;
		grayelecidleinferselout	:	OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		hipdatain	:	IN STD_LOGIC_VECTOR(9 DOWNTO 0) := (OTHERS => '0');
		hipdetectrxloop	:	IN STD_LOGIC := '0';
		hipelecidleinfersel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		hipforceelecidle	:	IN STD_LOGIC := '0';
		hippowerdn	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		hiptxclkout	:	OUT STD_LOGIC;
		invpol	:	IN STD_LOGIC := '0';
		localrefclk	:	IN STD_LOGIC := '0';
		parallelfdbkout	:	OUT STD_LOGIC_VECTOR(19 DOWNTO 0);
		phfifooverflow	:	OUT STD_LOGIC;
		phfiforddisable	:	IN STD_LOGIC := '0';
		phfiforddisableout	:	OUT STD_LOGIC;
		phfiforeset	:	IN STD_LOGIC := '0';
		phfiforesetout	:	OUT STD_LOGIC;
		phfifounderflow	:	OUT STD_LOGIC;
		phfifowrenable	:	IN STD_LOGIC := '1';
		phfifowrenableout	:	OUT STD_LOGIC;
		phfifox4bytesel	:	IN STD_LOGIC := '0';
		phfifox4rdclk	:	IN STD_LOGIC := '0';
		phfifox4rdenable	:	IN STD_LOGIC := '0';
		phfifox4wrenable	:	IN STD_LOGIC := '0';
		pipeenrevparallellpbkout	:	OUT STD_LOGIC;
		pipepowerdownout	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		pipepowerstateout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		pipestatetransdone	:	IN STD_LOGIC := '0';
		pipetxswing	:	IN STD_LOGIC := '0';
		powerdn	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		prbscidenable	:	IN STD_LOGIC := '0';
		quadreset	:	IN STD_LOGIC := '0';
		rdenablesync	:	OUT STD_LOGIC;
		refclk	:	IN STD_LOGIC := '0';
		revparallelfdbk	:	IN STD_LOGIC_VECTOR(19 DOWNTO 0) := (OTHERS => '0');
		txdetectrx	:	OUT STD_LOGIC;
		xgmctrl	:	IN STD_LOGIC := '0';
		xgmctrlenable	:	OUT STD_LOGIC;
		xgmdatain	:	IN STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		xgmdataout	:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  cycloneiv_hssi_tx_pma
	 GENERIC 
	 (
		channel_number	:	NATURAL := 0;
		common_mode	:	STRING := "0.65V";
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		effective_data_rate	:	STRING := "UNUSED";
		enable_diagnostic_loopback	:	STRING := "false";
		enable_reverse_serial_loopback	:	STRING := "false";
		enable_txclkout_loopback	:	STRING := "false";
		logical_channel_address	:	NATURAL := 0;
		preemp_tap_1	:	NATURAL := 0;
		protocol_hint	:	STRING := "basic";
		rx_detect	:	NATURAL := 0;
		serialization_factor	:	NATURAL := 8;
		slew_rate	:	STRING := "low";
		termination	:	STRING := "OCT 100 Ohms";
		use_external_termination	:	STRING := "false";
		use_rx_detect	:	STRING := "false";
		vod_selection	:	NATURAL := 0;
		lpm_type	:	STRING := "cycloneiv_hssi_tx_pma"
	 );
	 PORT
	 ( 
		cgbpowerdn	:	IN STD_LOGIC := '0';
		clockout	:	OUT STD_LOGIC;
		datain	:	IN STD_LOGIC_VECTOR(9 DOWNTO 0) := (OTHERS => '0');
		dataout	:	OUT STD_LOGIC;
		detectrxpowerdown	:	IN STD_LOGIC := '0';
		diagnosticlpbkin	:	IN STD_LOGIC := '0';
		dpriodisable	:	IN STD_LOGIC := '0';
		dprioin	:	IN STD_LOGIC_VECTOR(299 DOWNTO 0) := (OTHERS => '0');
		dprioout	:	OUT STD_LOGIC_VECTOR(299 DOWNTO 0);
		fastrefclk0in	:	IN STD_LOGIC := '0';
		forceelecidle	:	IN STD_LOGIC := '0';
		powerdn	:	IN STD_LOGIC := '0';
		refclk0in	:	IN STD_LOGIC := '0';
		refclk0inpulse	:	IN STD_LOGIC := '0';
		reverselpbkin	:	IN STD_LOGIC := '0';
		rxdetectclk	:	IN STD_LOGIC := '0';
		rxdetecten	:	IN STD_LOGIC := '0';
		rxdetectvalidout	:	OUT STD_LOGIC;
		rxfoundout	:	OUT STD_LOGIC;
		seriallpbkout	:	OUT STD_LOGIC;
		txpmareset	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	cal_blk_powerdown <= '0';
	cent_unit_quadresetout <= ( "000" & wire_cent_unit0_quadresetout);
	cent_unit_txdetectrxpowerdn <= ( wire_cent_unit0_txdetectrxpowerdown(3 DOWNTO 0));
	cent_unit_txdividerpowerdown <= ( wire_cent_unit0_txdividerpowerdown(3 DOWNTO 0));
	cent_unit_txobpowerdn <= ( wire_cent_unit0_txobpowerdown(3 DOWNTO 0));
	gxb_powerdown <= (OTHERS => '0');
	nonusertocmu_out(0) <= ( wire_cal_blk0_nonusertocmu);
	pll_locked(0) <= ( wire_pll0_locked);
	pll_powerdown <= (OTHERS => '0');
	reconfig_clk <= '0';
	tx_analogreset_out <= ( wire_cent_unit0_txanalogresetout(3 DOWNTO 0));
	tx_clkout <= ( tx_core_clkout_wire(3 DOWNTO 0));
	tx_clkout_int_wire <= ( wire_transmit_pcs3_clkout & wire_transmit_pcs2_clkout & wire_transmit_pcs1_clkout & wire_transmit_pcs0_clkout);
	tx_core_clkout_wire <= ( tx_clkout_int_wire(0) & tx_clkout_int_wire(0) & tx_clkout_int_wire(0) & tx_clkout_int_wire(0));
	tx_coreclk_in <= ( tx_clkout_int_wire(3 DOWNTO 0));
	tx_datain_wire <= ( tx_datain(63 DOWNTO 0));
	tx_dataout <= ( txdataout(3 DOWNTO 0));
	tx_dataout_pcs_to_pma <= ( wire_transmit_pcs3_dataout(9 DOWNTO 0) & wire_transmit_pcs2_dataout(9 DOWNTO 0) & wire_transmit_pcs1_dataout(9 DOWNTO 0) & wire_transmit_pcs0_dataout(9 DOWNTO 0));
	tx_digitalreset_in <= ( tx_digitalreset(3 DOWNTO 0));
	tx_digitalreset_out <= ( wire_cent_unit0_txdigitalresetout(3 DOWNTO 0));
	tx_forcedisp_wire <= ( "00" & "00" & "00" & "00");
	tx_invpolarity <= (OTHERS => '0');
	tx_localrefclk <= ( wire_transmit_pma3_clockout & wire_transmit_pma2_clockout & wire_transmit_pma1_clockout & wire_transmit_pma0_clockout);
	tx_phfiforeset <= (OTHERS => '0');
	tx_pma_fastrefclk0in <= ( wire_pll0_clk(0) & wire_pll0_clk(0) & wire_pll0_clk(0) & wire_pll0_clk(0));
	tx_pma_refclk0in <= ( wire_pll0_clk(1) & wire_pll0_clk(1) & wire_pll0_clk(1) & wire_pll0_clk(1));
	tx_pma_refclk0inpulse <= ( wire_pll0_clk(2) & wire_pll0_clk(2) & wire_pll0_clk(2) & wire_pll0_clk(2));
	tx_seriallpbkout <= ( wire_transmit_pma3_seriallpbkout & wire_transmit_pma2_seriallpbkout & wire_transmit_pma1_seriallpbkout & wire_transmit_pma0_seriallpbkout);
	txdataout <= ( wire_transmit_pma3_dataout & wire_transmit_pma2_dataout & wire_transmit_pma1_dataout & wire_transmit_pma0_dataout);
	txdetectrxout <= ( wire_transmit_pcs3_txdetectrx & wire_transmit_pcs2_txdetectrx & wire_transmit_pcs1_txdetectrx & wire_transmit_pcs0_txdetectrx);
	wire_pll0_areset <= wire_w_lg_w_pll_areset_range39w40w(0);
	wire_w_lg_w_pll_areset_range39w40w(0) <= pll_areset(0) OR pll_powerdown(0);
	wire_pll0_inclk <= ( "0" & pll_inclk(0));
	pll0 :  altpll
	  GENERIC MAP (
		bandwidth_type => "AUTO",
		clk0_divide_by => 5,
		clk0_multiply_by => 32,
		clk1_divide_by => 25,
		clk1_multiply_by => 32,
		clk2_divide_by => 25,
		clk2_duty_cycle => 20,
		clk2_multiply_by => 32,
		DPA_DIVIDE_BY => 5,
		DPA_MULTIPLY_BY => 32,
		inclk0_input_frequency => 10000,
		operation_mode => "no_compensation",
		INTENDED_DEVICE_FAMILY => "Cyclone IV GX"
	  )
	  PORT MAP ( 
		areset => wire_pll0_areset,
		clk => wire_pll0_clk,
		fref => wire_pll0_fref,
		icdrclk => wire_pll0_icdrclk,
		inclk => wire_pll0_inclk,
		locked => wire_pll0_locked
	  );
	cal_blk0 :  cycloneiv_hssi_calibration_block
	  PORT MAP ( 
		clk => cal_blk_clk,
		nonusertocmu => wire_cal_blk0_nonusertocmu,
		powerdn => cal_blk_powerdown
	  );
	wire_cent_unit0_adet <= (OTHERS => '0');
	wire_cent_unit0_rdalign <= (OTHERS => '0');
	wire_cent_unit0_rxctrl <= (OTHERS => '0');
	wire_cent_unit0_rxdatain <= (OTHERS => '0');
	wire_cent_unit0_rxdatavalid <= (OTHERS => '0');
	wire_cent_unit0_rxrunningdisp <= (OTHERS => '0');
	wire_cent_unit0_syncstatus <= (OTHERS => '0');
	wire_cent_unit0_txctrl <= (OTHERS => '0');
	wire_cent_unit0_txdatain <= (OTHERS => '0');
	wire_cent_unit0_txdigitalreset <= ( tx_digitalreset_in(3 DOWNTO 0));
	cent_unit0 :  cycloneiv_hssi_cmu
	  GENERIC MAP (
		auto_spd_deassert_ph_fifo_rst_count => 8,
		auto_spd_phystatus_notify_count => 14,
		devaddr => ((((starting_channel_number / 4) + 0) MOD 32) + 1),
		dprio_config_mode => "000000",
		in_xaui_mode => "false",
		portaddr => (((starting_channel_number + 0) / 128) + 1),
		rx0_ph_fifo_reg_mode => "false",
		tx0_channel_bonding => "none",
		tx0_rd_clk_mux_select => "central",
		tx0_reset_clock_output_during_digital_reset => "false",
		tx0_use_double_data_mode => "true",
		tx0_wr_clk_mux_select => "core_clk",
		use_coreclk_out_post_divider => "false",
		use_deskew_fifo => "false"
	  )
	  PORT MAP ( 
		adet => wire_cent_unit0_adet,
		dpclk => reconfig_clk,
		dpriodisable => wire_vcc,
		dprioin => wire_gnd,
		dprioload => wire_gnd,
		nonuserfromcal => nonusertocmu_out(0),
		quadreset => gxb_powerdown(0),
		quadresetout => wire_cent_unit0_quadresetout,
		rdalign => wire_cent_unit0_rdalign,
		rdenablesync => wire_gnd,
		recovclk => wire_gnd,
		rxctrl => wire_cent_unit0_rxctrl,
		rxdatain => wire_cent_unit0_rxdatain,
		rxdatavalid => wire_cent_unit0_rxdatavalid,
		rxrunningdisp => wire_cent_unit0_rxrunningdisp,
		syncstatus => wire_cent_unit0_syncstatus,
		txanalogresetout => wire_cent_unit0_txanalogresetout,
		txctrl => wire_cent_unit0_txctrl,
		txdatain => wire_cent_unit0_txdatain,
		txdetectrxpowerdown => wire_cent_unit0_txdetectrxpowerdown,
		txdigitalreset => wire_cent_unit0_txdigitalreset,
		txdigitalresetout => wire_cent_unit0_txdigitalresetout,
		txdividerpowerdown => wire_cent_unit0_txdividerpowerdown,
		txobpowerdown => wire_cent_unit0_txobpowerdown
	  );
	wire_transmit_pcs0_ctrlenable <= ( tx_ctrlenable(1 DOWNTO 0));
	wire_transmit_pcs0_datain <= ( "0000" & tx_datain_wire(15 DOWNTO 0));
	wire_transmit_pcs0_datainfull <= (OTHERS => '0');
	wire_transmit_pcs0_forcedisp <= ( tx_forcedisp_wire(1 DOWNTO 0));
	wire_transmit_pcs0_powerdn <= (OTHERS => '0');
	wire_transmit_pcs0_revparallelfdbk <= (OTHERS => '0');
	transmit_pcs0 :  cycloneiv_hssi_tx_pcs
	  GENERIC MAP (
		allow_polarity_inversion => "false",
		bitslip_enable => "false",
		channel_bonding => "none",
		channel_number => ((starting_channel_number + 0) MOD 4),
		channel_width => 16,
		core_clock_0ppm => "false",
		datapath_low_latency_mode => "false",
		datapath_protocol => "basic",
		disable_ph_low_latency_mode => "false",
		disparity_mode => "none",
		dprio_config_mode => "000000",
		elec_idle_delay => 6,
		enable_bit_reversal => "false",
		enable_idle_selection => "false",
		enable_reverse_parallel_loopback => "false",
		enable_self_test_mode => "false",
		enc_8b_10b_compatibility_mode => "true",
		enc_8b_10b_mode => "normal",
		hip_enable => "false",
		ph_fifo_reg_mode => "false",
		prbs_cid_pattern => "false",
		protocol_hint => "basic",
		refclk_select => "local",
		self_test_mode => "incremental",
		use_double_data_mode => "true",
		wr_clk_mux_select => "core_clk"
	  )
	  PORT MAP ( 
		clkout => wire_transmit_pcs0_clkout,
		coreclk => tx_coreclk_in(0),
		ctrlenable => wire_transmit_pcs0_ctrlenable,
		datain => wire_transmit_pcs0_datain,
		datainfull => wire_transmit_pcs0_datainfull,
		dataout => wire_transmit_pcs0_dataout,
		detectrxloop => wire_gnd,
		digitalreset => tx_digitalreset_out(0),
		dpriodisable => wire_vcc,
		enrevparallellpbk => wire_gnd,
		forcedisp => wire_transmit_pcs0_forcedisp,
		invpol => tx_invpolarity(0),
		localrefclk => tx_localrefclk(0),
		phfiforddisable => wire_gnd,
		phfiforeset => tx_phfiforeset(0),
		phfifowrenable => wire_vcc,
		pipestatetransdone => wire_gnd,
		powerdn => wire_transmit_pcs0_powerdn,
		quadreset => cent_unit_quadresetout(0),
		revparallelfdbk => wire_transmit_pcs0_revparallelfdbk,
		txdetectrx => wire_transmit_pcs0_txdetectrx
	  );
	wire_transmit_pcs1_ctrlenable <= ( tx_ctrlenable(3 DOWNTO 2));
	wire_transmit_pcs1_datain <= ( "0000" & tx_datain_wire(31 DOWNTO 16));
	wire_transmit_pcs1_datainfull <= (OTHERS => '0');
	wire_transmit_pcs1_forcedisp <= ( tx_forcedisp_wire(3 DOWNTO 2));
	wire_transmit_pcs1_powerdn <= (OTHERS => '0');
	wire_transmit_pcs1_revparallelfdbk <= (OTHERS => '0');
	transmit_pcs1 :  cycloneiv_hssi_tx_pcs
	  GENERIC MAP (
		allow_polarity_inversion => "false",
		bitslip_enable => "false",
		channel_bonding => "none",
		channel_number => ((starting_channel_number + 1) MOD 4),
		channel_width => 16,
		core_clock_0ppm => "false",
		datapath_low_latency_mode => "false",
		datapath_protocol => "basic",
		disable_ph_low_latency_mode => "false",
		disparity_mode => "none",
		dprio_config_mode => "000000",
		elec_idle_delay => 6,
		enable_bit_reversal => "false",
		enable_idle_selection => "false",
		enable_reverse_parallel_loopback => "false",
		enable_self_test_mode => "false",
		enc_8b_10b_compatibility_mode => "true",
		enc_8b_10b_mode => "normal",
		hip_enable => "false",
		ph_fifo_reg_mode => "false",
		prbs_cid_pattern => "false",
		protocol_hint => "basic",
		refclk_select => "local",
		self_test_mode => "incremental",
		use_double_data_mode => "true",
		wr_clk_mux_select => "core_clk"
	  )
	  PORT MAP ( 
		clkout => wire_transmit_pcs1_clkout,
		coreclk => tx_coreclk_in(1),
		ctrlenable => wire_transmit_pcs1_ctrlenable,
		datain => wire_transmit_pcs1_datain,
		datainfull => wire_transmit_pcs1_datainfull,
		dataout => wire_transmit_pcs1_dataout,
		detectrxloop => wire_gnd,
		digitalreset => tx_digitalreset_out(1),
		dpriodisable => wire_vcc,
		enrevparallellpbk => wire_gnd,
		forcedisp => wire_transmit_pcs1_forcedisp,
		invpol => tx_invpolarity(1),
		localrefclk => tx_localrefclk(1),
		phfiforddisable => wire_gnd,
		phfiforeset => tx_phfiforeset(1),
		phfifowrenable => wire_vcc,
		pipestatetransdone => wire_gnd,
		powerdn => wire_transmit_pcs1_powerdn,
		quadreset => cent_unit_quadresetout(0),
		revparallelfdbk => wire_transmit_pcs1_revparallelfdbk,
		txdetectrx => wire_transmit_pcs1_txdetectrx
	  );
	wire_transmit_pcs2_ctrlenable <= ( tx_ctrlenable(5 DOWNTO 4));
	wire_transmit_pcs2_datain <= ( "0000" & tx_datain_wire(47 DOWNTO 32));
	wire_transmit_pcs2_datainfull <= (OTHERS => '0');
	wire_transmit_pcs2_forcedisp <= ( tx_forcedisp_wire(5 DOWNTO 4));
	wire_transmit_pcs2_powerdn <= (OTHERS => '0');
	wire_transmit_pcs2_revparallelfdbk <= (OTHERS => '0');
	transmit_pcs2 :  cycloneiv_hssi_tx_pcs
	  GENERIC MAP (
		allow_polarity_inversion => "false",
		bitslip_enable => "false",
		channel_bonding => "none",
		channel_number => ((starting_channel_number + 2) MOD 4),
		channel_width => 16,
		core_clock_0ppm => "false",
		datapath_low_latency_mode => "false",
		datapath_protocol => "basic",
		disable_ph_low_latency_mode => "false",
		disparity_mode => "none",
		dprio_config_mode => "000000",
		elec_idle_delay => 6,
		enable_bit_reversal => "false",
		enable_idle_selection => "false",
		enable_reverse_parallel_loopback => "false",
		enable_self_test_mode => "false",
		enc_8b_10b_compatibility_mode => "true",
		enc_8b_10b_mode => "normal",
		hip_enable => "false",
		ph_fifo_reg_mode => "false",
		prbs_cid_pattern => "false",
		protocol_hint => "basic",
		refclk_select => "local",
		self_test_mode => "incremental",
		use_double_data_mode => "true",
		wr_clk_mux_select => "core_clk"
	  )
	  PORT MAP ( 
		clkout => wire_transmit_pcs2_clkout,
		coreclk => tx_coreclk_in(2),
		ctrlenable => wire_transmit_pcs2_ctrlenable,
		datain => wire_transmit_pcs2_datain,
		datainfull => wire_transmit_pcs2_datainfull,
		dataout => wire_transmit_pcs2_dataout,
		detectrxloop => wire_gnd,
		digitalreset => tx_digitalreset_out(2),
		dpriodisable => wire_vcc,
		enrevparallellpbk => wire_gnd,
		forcedisp => wire_transmit_pcs2_forcedisp,
		invpol => tx_invpolarity(2),
		localrefclk => tx_localrefclk(2),
		phfiforddisable => wire_gnd,
		phfiforeset => tx_phfiforeset(2),
		phfifowrenable => wire_vcc,
		pipestatetransdone => wire_gnd,
		powerdn => wire_transmit_pcs2_powerdn,
		quadreset => cent_unit_quadresetout(0),
		revparallelfdbk => wire_transmit_pcs2_revparallelfdbk,
		txdetectrx => wire_transmit_pcs2_txdetectrx
	  );
	wire_transmit_pcs3_ctrlenable <= ( tx_ctrlenable(7 DOWNTO 6));
	wire_transmit_pcs3_datain <= ( "0000" & tx_datain_wire(63 DOWNTO 48));
	wire_transmit_pcs3_datainfull <= (OTHERS => '0');
	wire_transmit_pcs3_forcedisp <= ( tx_forcedisp_wire(7 DOWNTO 6));
	wire_transmit_pcs3_powerdn <= (OTHERS => '0');
	wire_transmit_pcs3_revparallelfdbk <= (OTHERS => '0');
	transmit_pcs3 :  cycloneiv_hssi_tx_pcs
	  GENERIC MAP (
		allow_polarity_inversion => "false",
		bitslip_enable => "false",
		channel_bonding => "none",
		channel_number => ((starting_channel_number + 3) MOD 4),
		channel_width => 16,
		core_clock_0ppm => "false",
		datapath_low_latency_mode => "false",
		datapath_protocol => "basic",
		disable_ph_low_latency_mode => "false",
		disparity_mode => "none",
		dprio_config_mode => "000000",
		elec_idle_delay => 6,
		enable_bit_reversal => "false",
		enable_idle_selection => "false",
		enable_reverse_parallel_loopback => "false",
		enable_self_test_mode => "false",
		enc_8b_10b_compatibility_mode => "true",
		enc_8b_10b_mode => "normal",
		hip_enable => "false",
		ph_fifo_reg_mode => "false",
		prbs_cid_pattern => "false",
		protocol_hint => "basic",
		refclk_select => "local",
		self_test_mode => "incremental",
		use_double_data_mode => "true",
		wr_clk_mux_select => "core_clk"
	  )
	  PORT MAP ( 
		clkout => wire_transmit_pcs3_clkout,
		coreclk => tx_coreclk_in(3),
		ctrlenable => wire_transmit_pcs3_ctrlenable,
		datain => wire_transmit_pcs3_datain,
		datainfull => wire_transmit_pcs3_datainfull,
		dataout => wire_transmit_pcs3_dataout,
		detectrxloop => wire_gnd,
		digitalreset => tx_digitalreset_out(3),
		dpriodisable => wire_vcc,
		enrevparallellpbk => wire_gnd,
		forcedisp => wire_transmit_pcs3_forcedisp,
		invpol => tx_invpolarity(3),
		localrefclk => tx_localrefclk(3),
		phfiforddisable => wire_gnd,
		phfiforeset => tx_phfiforeset(3),
		phfifowrenable => wire_vcc,
		pipestatetransdone => wire_gnd,
		powerdn => wire_transmit_pcs3_powerdn,
		quadreset => cent_unit_quadresetout(0),
		revparallelfdbk => wire_transmit_pcs3_revparallelfdbk,
		txdetectrx => wire_transmit_pcs3_txdetectrx
	  );
	wire_transmit_pma0_datain <= ( tx_dataout_pcs_to_pma(9 DOWNTO 0));
	transmit_pma0 :  cycloneiv_hssi_tx_pma
	  GENERIC MAP (
		channel_number => ((starting_channel_number + 0) MOD 4),
		common_mode => "0.65V",
		dprio_config_mode => "000000",
		effective_data_rate => "1280 Mbps",
		enable_diagnostic_loopback => "false",
		enable_reverse_serial_loopback => "false",
		logical_channel_address => (starting_channel_number + 0),
		preemp_tap_1 => 0,
		protocol_hint => "basic",
		rx_detect => 0,
		serialization_factor => 10,
		slew_rate => "low",
		termination => "OCT 100 Ohms",
		use_external_termination => "false",
		use_rx_detect => "false",
		vod_selection => 6
	  )
	  PORT MAP ( 
		cgbpowerdn => cent_unit_txdividerpowerdown(0),
		clockout => wire_transmit_pma0_clockout,
		datain => wire_transmit_pma0_datain,
		dataout => wire_transmit_pma0_dataout,
		detectrxpowerdown => cent_unit_txdetectrxpowerdn(0),
		diagnosticlpbkin => tx_diagnosticlpbkin(0),
		dpriodisable => wire_vcc,
		fastrefclk0in => tx_pma_fastrefclk0in(0),
		forceelecidle => wire_gnd,
		powerdn => cent_unit_txobpowerdn(0),
		refclk0in => tx_pma_refclk0in(0),
		refclk0inpulse => tx_pma_refclk0inpulse(0),
		rxdetecten => txdetectrxout(0),
		seriallpbkout => wire_transmit_pma0_seriallpbkout,
		txpmareset => tx_analogreset_out(0)
	  );
	wire_transmit_pma1_datain <= ( tx_dataout_pcs_to_pma(19 DOWNTO 10));
	transmit_pma1 :  cycloneiv_hssi_tx_pma
	  GENERIC MAP (
		channel_number => ((starting_channel_number + 1) MOD 4),
		common_mode => "0.65V",
		dprio_config_mode => "000000",
		effective_data_rate => "1280 Mbps",
		enable_diagnostic_loopback => "false",
		enable_reverse_serial_loopback => "false",
		logical_channel_address => (starting_channel_number + 1),
		preemp_tap_1 => 0,
		protocol_hint => "basic",
		rx_detect => 0,
		serialization_factor => 10,
		slew_rate => "low",
		termination => "OCT 100 Ohms",
		use_external_termination => "false",
		use_rx_detect => "false",
		vod_selection => 6
	  )
	  PORT MAP ( 
		cgbpowerdn => cent_unit_txdividerpowerdown(1),
		clockout => wire_transmit_pma1_clockout,
		datain => wire_transmit_pma1_datain,
		dataout => wire_transmit_pma1_dataout,
		detectrxpowerdown => cent_unit_txdetectrxpowerdn(1),
		diagnosticlpbkin => tx_diagnosticlpbkin(1),
		dpriodisable => wire_vcc,
		fastrefclk0in => tx_pma_fastrefclk0in(1),
		forceelecidle => wire_gnd,
		powerdn => cent_unit_txobpowerdn(1),
		refclk0in => tx_pma_refclk0in(1),
		refclk0inpulse => tx_pma_refclk0inpulse(1),
		rxdetecten => txdetectrxout(1),
		seriallpbkout => wire_transmit_pma1_seriallpbkout,
		txpmareset => tx_analogreset_out(1)
	  );
	wire_transmit_pma2_datain <= ( tx_dataout_pcs_to_pma(29 DOWNTO 20));
	transmit_pma2 :  cycloneiv_hssi_tx_pma
	  GENERIC MAP (
		channel_number => ((starting_channel_number + 2) MOD 4),
		common_mode => "0.65V",
		dprio_config_mode => "000000",
		effective_data_rate => "1280 Mbps",
		enable_diagnostic_loopback => "false",
		enable_reverse_serial_loopback => "false",
		logical_channel_address => (starting_channel_number + 2),
		preemp_tap_1 => 0,
		protocol_hint => "basic",
		rx_detect => 0,
		serialization_factor => 10,
		slew_rate => "low",
		termination => "OCT 100 Ohms",
		use_external_termination => "false",
		use_rx_detect => "false",
		vod_selection => 6
	  )
	  PORT MAP ( 
		cgbpowerdn => cent_unit_txdividerpowerdown(2),
		clockout => wire_transmit_pma2_clockout,
		datain => wire_transmit_pma2_datain,
		dataout => wire_transmit_pma2_dataout,
		detectrxpowerdown => cent_unit_txdetectrxpowerdn(2),
		diagnosticlpbkin => tx_diagnosticlpbkin(2),
		dpriodisable => wire_vcc,
		fastrefclk0in => tx_pma_fastrefclk0in(2),
		forceelecidle => wire_gnd,
		powerdn => cent_unit_txobpowerdn(2),
		refclk0in => tx_pma_refclk0in(2),
		refclk0inpulse => tx_pma_refclk0inpulse(2),
		rxdetecten => txdetectrxout(2),
		seriallpbkout => wire_transmit_pma2_seriallpbkout,
		txpmareset => tx_analogreset_out(2)
	  );
	wire_transmit_pma3_datain <= ( tx_dataout_pcs_to_pma(39 DOWNTO 30));
	transmit_pma3 :  cycloneiv_hssi_tx_pma
	  GENERIC MAP (
		channel_number => ((starting_channel_number + 3) MOD 4),
		common_mode => "0.65V",
		dprio_config_mode => "000000",
		effective_data_rate => "1280 Mbps",
		enable_diagnostic_loopback => "false",
		enable_reverse_serial_loopback => "false",
		logical_channel_address => (starting_channel_number + 3),
		preemp_tap_1 => 0,
		protocol_hint => "basic",
		rx_detect => 0,
		serialization_factor => 10,
		slew_rate => "low",
		termination => "OCT 100 Ohms",
		use_external_termination => "false",
		use_rx_detect => "false",
		vod_selection => 6
	  )
	  PORT MAP ( 
		cgbpowerdn => cent_unit_txdividerpowerdown(3),
		clockout => wire_transmit_pma3_clockout,
		datain => wire_transmit_pma3_datain,
		dataout => wire_transmit_pma3_dataout,
		detectrxpowerdown => cent_unit_txdetectrxpowerdn(3),
		diagnosticlpbkin => tx_diagnosticlpbkin(3),
		dpriodisable => wire_vcc,
		fastrefclk0in => tx_pma_fastrefclk0in(3),
		forceelecidle => wire_gnd,
		powerdn => cent_unit_txobpowerdn(3),
		refclk0in => tx_pma_refclk0in(3),
		refclk0inpulse => tx_pma_refclk0inpulse(3),
		rxdetecten => txdetectrxout(3),
		seriallpbkout => wire_transmit_pma3_seriallpbkout,
		txpmareset => tx_analogreset_out(3)
	  );

 END RTL; --ALTGX_TX_alt_c3gxb
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ALTGX_TX IS
	PORT
	(
		cal_blk_clk		: IN STD_LOGIC ;
		pll_areset		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		pll_inclk		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		tx_ctrlenable		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		tx_datain		: IN STD_LOGIC_VECTOR (63 DOWNTO 0);
		tx_digitalreset		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		pll_locked		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		tx_clkout		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		tx_dataout		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
END ALTGX_TX;


ARCHITECTURE RTL OF altgx_tx IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (3 DOWNTO 0);



	COMPONENT ALTGX_TX_alt_c3gxb
	PORT (
			cal_blk_clk	: IN STD_LOGIC ;
			pll_areset	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			pll_inclk	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			tx_ctrlenable	: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			tx_datain	: IN STD_LOGIC_VECTOR (63 DOWNTO 0);
			tx_digitalreset	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			pll_locked	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			tx_clkout	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			tx_dataout	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	pll_locked    <= sub_wire0(0 DOWNTO 0);
	tx_clkout    <= sub_wire1(3 DOWNTO 0);
	tx_dataout    <= sub_wire2(3 DOWNTO 0);

	ALTGX_TX_alt_c3gxb_component : ALTGX_TX_alt_c3gxb
	PORT MAP (
		cal_blk_clk => cal_blk_clk,
		pll_areset => pll_areset,
		pll_inclk => pll_inclk,
		tx_ctrlenable => tx_ctrlenable,
		tx_datain => tx_datain,
		tx_digitalreset => tx_digitalreset,
		pll_locked => sub_wire0,
		tx_clkout => sub_wire1,
		tx_dataout => sub_wire2
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: PRIVATE: NUM_KEYS NUMERIC "0"
-- Retrieval info: PRIVATE: RECONFIG_PROTOCOL STRING "BASIC"
-- Retrieval info: PRIVATE: RECONFIG_SUBPROTOCOL STRING "none"
-- Retrieval info: PRIVATE: RX_ENABLE_DC_COUPLING STRING "false"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE STRING "1280"
-- Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE_ENABLE STRING "0"
-- Retrieval info: PRIVATE: WIZ_DATA_RATE STRING "1280"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INCLK_FREQ_ARRAY STRING "100"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A STRING "2000"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A_UNIT STRING "Mbps"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B STRING "100"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B_UNIT STRING "MHz"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_SELECTION NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_FREQ STRING "50.526315"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_ENABLE_EQUALIZER_CTRL NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_EQUALIZER_CTRL_SETTING NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_FORCE_DEFAULT_SETTINGS NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_INCLK_FREQ STRING "100.0"
-- Retrieval info: PRIVATE: WIZ_INCLK_FREQ_ARRAY STRING "50.526315 51.2 51.891891 53.333333 54.857142 55.652173 56.470588 58.181818 60.0 60.95238 61.935483 64.0 65.641025 66.206896 67.368421 68.571428 69.189189 71.111111 73.142857 73.846153"
-- Retrieval info: PRIVATE: WIZ_INPUT_A STRING "1280"
-- Retrieval info: PRIVATE: WIZ_INPUT_A_UNIT STRING "Mbps"
-- Retrieval info: PRIVATE: WIZ_INPUT_B STRING "100.0"
-- Retrieval info: PRIVATE: WIZ_INPUT_B_UNIT STRING "MHz"
-- Retrieval info: PRIVATE: WIZ_INPUT_SELECTION NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_SUBPROTOCOL STRING "None"
-- Retrieval info: PRIVATE: WIZ_WORD_ALIGN_FLIP_PATTERN STRING "0"
-- Retrieval info: CONSTANT: EFFECTIVE_DATA_RATE STRING "1280 Mbps"
-- Retrieval info: CONSTANT: ENABLE_LC_TX_PLL STRING "false"
-- Retrieval info: CONSTANT: ENABLE_PLL_INCLK_ALT_DRIVE_RX_CRU STRING "true"
-- Retrieval info: CONSTANT: ENABLE_PLL_INCLK_DRIVE_RX_CRU STRING "true"
-- Retrieval info: CONSTANT: GX_CHANNEL_TYPE STRING ""
-- Retrieval info: CONSTANT: INPUT_CLOCK_FREQUENCY STRING "100.0 MHz"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_SPEED_GRADE STRING "6"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_VARIANT STRING "ANY"
-- Retrieval info: CONSTANT: LOOPBACK_MODE STRING "none"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "alt_c3gxb"
-- Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "4"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "tx"
-- Retrieval info: CONSTANT: PLL_BANDWIDTH_TYPE STRING "Auto"
-- Retrieval info: CONSTANT: PLL_CONTROL_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: PLL_INCLK_PERIOD NUMERIC "10000"
-- Retrieval info: CONSTANT: PLL_PFD_FB_MODE STRING "internal"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_1STPOSTTAP_SETTING NUMERIC "0"
-- Retrieval info: CONSTANT: PROTOCOL STRING "basic"
-- Retrieval info: CONSTANT: RECONFIG_DPRIO_MODE NUMERIC "0"
-- Retrieval info: CONSTANT: RX_CRU_INCLOCK0_PERIOD NUMERIC "10000"
-- Retrieval info: CONSTANT: TRANSMITTER_TERMINATION STRING "oct_100_ohms"
-- Retrieval info: CONSTANT: TX_8B_10B_MODE STRING "normal"
-- Retrieval info: CONSTANT: TX_ALLOW_POLARITY_INVERSION STRING "false"
-- Retrieval info: CONSTANT: TX_CHANNEL_WIDTH NUMERIC "16"
-- Retrieval info: CONSTANT: TX_CLKOUT_WIDTH NUMERIC "4"
-- Retrieval info: CONSTANT: TX_COMMON_MODE STRING "0.65v"
-- Retrieval info: CONSTANT: TX_DATAPATH_LOW_LATENCY_MODE STRING "false"
-- Retrieval info: CONSTANT: TX_DATA_RATE NUMERIC "1280"
-- Retrieval info: CONSTANT: TX_DATA_RATE_REMAINDER NUMERIC "0"
-- Retrieval info: CONSTANT: TX_DIGITALRESET_PORT_WIDTH NUMERIC "4"
-- Retrieval info: CONSTANT: TX_ENABLE_BIT_REVERSAL STRING "false"
-- Retrieval info: CONSTANT: TX_ENABLE_SELF_TEST_MODE STRING "false"
-- Retrieval info: CONSTANT: TX_FLIP_TX_IN STRING "false"
-- Retrieval info: CONSTANT: TX_FORCE_DISPARITY_MODE STRING "false"
-- Retrieval info: CONSTANT: TX_PLL_BANDWIDTH_TYPE STRING "Auto"
-- Retrieval info: CONSTANT: TX_PLL_INCLK0_PERIOD NUMERIC "10000"
-- Retrieval info: CONSTANT: TX_PLL_TYPE STRING "CMU"
-- Retrieval info: CONSTANT: TX_SLEW_RATE STRING "low"
-- Retrieval info: CONSTANT: TX_TRANSMIT_PROTOCOL STRING "basic"
-- Retrieval info: CONSTANT: TX_USE_CORECLK STRING "false"
-- Retrieval info: CONSTANT: TX_USE_DOUBLE_DATA_MODE STRING "true"
-- Retrieval info: CONSTANT: TX_USE_SERIALIZER_DOUBLE_DATA_MODE STRING "false"
-- Retrieval info: CONSTANT: USE_CALIBRATION_BLOCK STRING "true"
-- Retrieval info: CONSTANT: VOD_CTRL_SETTING NUMERIC "6"
-- Retrieval info: CONSTANT: gxb_powerdown_width NUMERIC "1"
-- Retrieval info: CONSTANT: iqtxrxclk_allowed STRING ""
-- Retrieval info: CONSTANT: number_of_quads NUMERIC "1"
-- Retrieval info: CONSTANT: pll_divide_by STRING "5"
-- Retrieval info: CONSTANT: pll_multiply_by STRING "32"
-- Retrieval info: CONSTANT: rx_enable_second_order_loop STRING "false"
-- Retrieval info: CONSTANT: rx_loop_1_digital_filter NUMERIC "8"
-- Retrieval info: CONSTANT: tx_bitslip_enable STRING "FALSE"
-- Retrieval info: CONSTANT: tx_dwidth_factor NUMERIC "2"
-- Retrieval info: CONSTANT: tx_use_external_termination STRING "false"
-- Retrieval info: USED_PORT: cal_blk_clk 0 0 0 0 INPUT NODEFVAL "cal_blk_clk"
-- Retrieval info: USED_PORT: pll_areset 0 0 1 0 INPUT NODEFVAL "pll_areset[0..0]"
-- Retrieval info: USED_PORT: pll_inclk 0 0 1 0 INPUT NODEFVAL "pll_inclk[0..0]"
-- Retrieval info: USED_PORT: pll_locked 0 0 1 0 OUTPUT NODEFVAL "pll_locked[0..0]"
-- Retrieval info: USED_PORT: tx_clkout 0 0 4 0 OUTPUT NODEFVAL "tx_clkout[3..0]"
-- Retrieval info: USED_PORT: tx_ctrlenable 0 0 8 0 INPUT NODEFVAL "tx_ctrlenable[7..0]"
-- Retrieval info: USED_PORT: tx_datain 0 0 64 0 INPUT NODEFVAL "tx_datain[63..0]"
-- Retrieval info: USED_PORT: tx_dataout 0 0 4 0 OUTPUT NODEFVAL "tx_dataout[3..0]"
-- Retrieval info: USED_PORT: tx_digitalreset 0 0 4 0 INPUT NODEFVAL "tx_digitalreset[3..0]"
-- Retrieval info: CONNECT: @cal_blk_clk 0 0 0 0 cal_blk_clk 0 0 0 0
-- Retrieval info: CONNECT: @pll_areset 0 0 1 0 pll_areset 0 0 1 0
-- Retrieval info: CONNECT: @pll_inclk 0 0 1 0 pll_inclk 0 0 1 0
-- Retrieval info: CONNECT: @tx_ctrlenable 0 0 8 0 tx_ctrlenable 0 0 8 0
-- Retrieval info: CONNECT: @tx_datain 0 0 64 0 tx_datain 0 0 64 0
-- Retrieval info: CONNECT: @tx_digitalreset 0 0 4 0 tx_digitalreset 0 0 4 0
-- Retrieval info: CONNECT: pll_locked 0 0 1 0 @pll_locked 0 0 1 0
-- Retrieval info: CONNECT: tx_clkout 0 0 4 0 @tx_clkout 0 0 4 0
-- Retrieval info: CONNECT: tx_dataout 0 0 4 0 @tx_dataout 0 0 4 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL ALTGX_TX.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ALTGX_TX.ppf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ALTGX_TX.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ALTGX_TX.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ALTGX_TX.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ALTGX_TX_inst.vhd FALSE
-- Retrieval info: CBX_MODULE_PREFIX: ON
