// Copyright (C) 1991-2014 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1.4
// ALTERA_TIMESTAMP:Thu Mar 13 15:23:43 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jxBhLqQfl3I+ugtXsiMbj9Bzg4qjCbQmu78wdON5kExMYww9vKR8uZ20UMbbYR6w
o3YPdnjHNLw62BXYDHuSFCl+R6t2qd0etcvUaHc47mfQka8qgvQiyCA3Bcc7MdoL
HYzhtBMuApmiGc9V3yovh/6wFQsD/qiLLF6MTj5gPl0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9664)
pqonU//ZayNgh1JJPEyetoxNk3ARG77y5foHY7yOnExiaIeWevcL+qJIKocksVTj
sELj7eXTqGdXMwou7VW7u6mpO+M5VLKNDIgRLMxXbPhTep8QlYR0KynO0FsuHG0/
9TT/nOkQnxTCZLvezweoKV2Ptp0dlf0GST3yKRc+0iIrsZYrhI2LtvcEyzzlKHHK
/Ib9JeG1+5Gp4gauY9QqevHQ/KphBNJ6LyAYBIuknS7VqFd+vcOAhRJg9XZq22OV
2eexkaVq/x1iFrXFQY2dod4DfQ6oCDXsq6le5j+JE85oIjjnAvAXr1m7NqdGWP7c
aoonIj3XShFuRLGtlWxfMZdv0EAStIbpRH2/JlzdnClEd0/LpUwiRK2vrEZVAnBM
JC0ZQ16QElenPHB2GwE9JNtDmxr9Nv2wnD0WkL50CjnHX7EkmVfqtOW9fPx5HlFp
XSRudt9SCmtxjVxZKEhjSW27HsLW8hQb1Xw9ZydystVlwgBDyu/wD/kCGC9vMQtp
iCCBMRzHmQc93wGOtssXjFirupi/3uO9EoANJODWDHgH0ugRAe7zzk4zgQg5i0ms
FH5DLdnV3qEXCZq3S/I0+96FGxbf8tpRQaeM1fRfghVeRzExWrO5rbvWdlYWuqHI
Ile6EY3i3lG57EK9qfMjgYxaQlX/+HjB8YZfuFLFfxyvIVztYLCqeCCdKYv4T8KD
WrGx+N4k4Hj99ZhXS/IJc1RnpjaJFTx+sAY3KAZsk5o8q/OaMY54bd1C9vUtA2+M
C2wjInW850PsrDnSAN2QN5s4qD3sia3VChas/MJI/RICVqVqoaPo7EGcUtcS/2Mu
q2tZ8poV4XnOOX44gJ/jZR63NcAk5dJzk6QiJYQzCdOAYvyYqqymVR8UQVeMHp6s
bHgrhKAKwUpMYOt5+T92EofldBqnkeKPziF7dQizoUrdLipxtO3OBJ+k+TC1l27w
MODKH8PakWwiVZKtqKqqESW8zX+5rNkmCn5xiMH6ZkiJ74av1asJMQuzMzA7SBnV
o6vbHHkruzv9wkHW/bkiHjztFJuzxQpbWZQ68vQHo7V7k04TjrDGm+UYX/3C+2la
5qZDkVoz9mTbiMfaEBkefaYHEfizm/6e1UZbsNy57yOrprCKuQX8H14aNu1YswKx
Ew1pjOkXICtxJyg2FZMPScNDIFCKXOyIdXxRsHoKsaYhu+Zfv15C3RGIUyvTg/Wu
pdyknE9HGuKdtHxcY/cB8w4+PF7GJZ5V03mibaKP6F3wzaZXCTxDg9YlDRbvffQA
Slx+UpJ6QSJbVtKcudDWpLbjJXukCXkndpfdx7E+2LP3CIfV+XNOUGG/Q8M8xehd
vv4kZK23SnEyKSBm+0SS4I3HpHEkEmPrbpsUJB6FRecXT4emLO4dndLrBhU19ec4
BPBL4fy7E5Z0c0Af7m6KOhW0/HVMsxXM0T/oVoHnv/2EdOT92Y1rpUogxnVRlPLa
25GCLD5BGzDHTSpJ8o5kQU/I4cMv+VDM3dMbywO6Lvwdavxj/cvDAaqev9MTXFG6
JsLowFZ65wvRRzCGqnQePZoMF6FMoVVYcNgpv45Qa3DKvQotb/nVzIk0D/7v8coM
xVG3ZkehT4faM/fdIo2iQe2Djtbe179ZRbz6Jw2lZDFc1hZZuJHGIFPszjRyuHAD
TKeKLIrn8K+1ocE4B2hJySSW1lfu/3B177iKq4RImenk0jCTmROOINodphAbY+Nn
t3AXgoCMsWqXllRhu9EYxpFuUYHDgMFw+OfanrBAxbDeSylGmKYwZNEEYdNz7KT+
/Rqgey4y+j7/pmdc41qL9F69sSeUCy49gL4h98aRvFCdO7uurP7e++HWj8KmJF/9
BjGzzB91CindxbZwIRm8mpNBNQGT2bYeS5Q7gikdttvbt5XxznmDgmVx+IG4DgCJ
HhRQMLrvJCCTs6nJJFzOJ7MSklPnnOmjmtz3RyZ2K5KIRH6c0t4Dd+zni3fe/ijB
kW0ks46XBQtGCJ6JCVbJTYb0STtnTeDfy6zoxi3BCfaa6Z3+dsUUDvJT1mRKiGJM
yFkAFp5fcox1rIJn103QXJu8qf3VCi5N2RfpIlmUcs00Z8IQ+GSciuneSpQw1Ds/
aF2QjYOBDel2xEDcN2CTKqR0Y2ehs6KHumKz8QbwP9ziYiqX8Jw/nsty/cS48QdE
udkVt6G7jm5gKvGHrxRkkrlh5DZIwtuMw++Wlp40xPu14HUDh/rXLy+GtYmsvL0Y
ddrg3ozc6w2l822wXmf2bBfG3iooe2NteRaoYUuvxiamcY0YmiXE0JfGxdFawAIn
5/MBza3pE6ozDqCI28ON19kHxbcUVdbjC34itQTkYEj7OiKoPG4aShvIPAs2ykjI
mMJbKCb42D1EpVVOF04CEU/e28HE86ly6GjhG6gky/OuinEPFbCpenGrkEdHf4KX
ZblQyZdz0gRuwUmy1EASYV43jLVYU7irTbdx6K5Z73yj9MvA2U18u1s4aGVWp5wO
0KehpWBJ2fdgIm5sVohvyO9n+CFRMImrOkeLE3ZCZW551hQH6vF0icYsCqgl+P6Y
aaogNLo84cBrRUHsF1EY9U2kBF952Hxu30JI1QDp/MouVkl2ORmZGhbONm5WP71s
/lDzZjVoIRtaEaPjzC5pZsDUMktEv3jN8/HAS0l3FVdFgvX35wlydE1mVzNoddmZ
4+KyCDwqdUwmoJRBkd+hRT6tP42Z1/Y6xcbY9teL54TVP0+Gx3U3g1Wa6E7YYl5N
zS+pcUNpc7DvkJB6P2LQvNtYE1qB602v/G2W2VTuzfygHNvnllTUGaIG12NKB9Ea
i8BxjHCeDF4KCAzRGZIlv5MXX+p2OB9OmWBxXyF4WNUE6udDP7LO1FE9NSFC8ApG
TAKoixMzIx83W1beAC/QQTRmV4M9N2SDpABrzV1si1dfdQZiNHgaoF57J92cOCTV
VNoBszvY2xSxMc2vC8YHCvYEmtfdRMZJDUmH/o0Sn4QDND7RDD10UqbwjEDrT6mS
wRH4cN4jKd42NNqNaRUlQ6GOiM706ewws9ZB61eOrQRXGHWAUwc9ecJlZKxZNaII
OkkatYuTleCmqEdQp9LVDMq+2Gh5YoKmHTiORSNMf0jDTb7vlJZE8ysOPmLlWEvS
idPRCiIdqL0L2JmgoT6gwKNwhWMqrgWclDGw92UvYPHJMWv/n8FY0SVrh5YQUyY3
mBa/QrXDU154jSsc9VVoWiVWyKrCqqVsijt4tivE/c1aEGu8tgWfGCL5f1NHNruD
koKq4F+xItBTEaQqTRcssibaIvSelu/S3qxixp9/Kqh/cZehXfhe9nOA6MNxp1e6
JxcoVNjXeQR92en6HnGfbARD192LMIMTjpRd+KC3fbPhEWnU05xSjKD+BZlghAzY
bYT6MM9oX2/yFTvV1HFuYGVcSCCT5QSRnCUQ6UzeEpOMr+2A0d37vYY9twq8D+zL
kSZ8lqTWInZI5dp0DDt9cpEw0DVD5aW+q2lFDbLUMv76pnaC5/i2cSn1Ai25Ojkf
RSsyYQIOq+s7IfmfB3HxoZv8bNkox5GSjeXCZljLYxlTgPlXe7vEimucl6WHoYa1
dlwuMHYpHBYj1ZmT+XpfIKRmhXEGkFsTRHgc/48/C5PFddSGoGjpZq6MpjRh9hp7
DIno8FhdnN7LqIbmgpp8tEc8st1kXJvqBCvi1fjzW0irHqh/PvIpU1aFmW40b+Kf
0al+ibbQbbhGdZmpto+j2E7dSij7c410rluL0lhCs1T6ek7c/iZUwgvL8w51HFsB
euWkyGYKHY7TEA0KC3Wnj2hqP4zj2KY3nIlsLRNZLFo3NJZI9sgRXbHVZbLy8RHB
FpokVhBHgKFJCbyuquJqMKJBnxsZWef8yffIV1kW8+tHFeKw6bEN/GMR/riHgUOX
DxgLPhk/ypmrtGPEGzpn91XmGDZ7CHL8PJc7kZksKgmIAjgJ/J7m+c9Fy1p0zO5C
GdoV04rLbKjgWx8BqTapMV8hz1Xf9+H8HQ03skb9jPlACajoKBvkzWQ+PM+YuEb9
lmvMBuX1ww9sVkcK0bngKvX6ux0euvIST/tQePJogw0nI663BfDH/A4zp226yxAa
/h/byCbeWJq3xoNr/oirEB7Y4Ny3UPfcOHY5hswjHEObhjPR3kN9IIfHGrk4eGwv
KJ4KO9auLpxLzvT/GPoFoYy5Wl8L3iCnHolhqYjLM6zyGu7X4pQXSJslrImAERTS
9eTqNdv+NgK296eHhEZnRVVobwZ2NRlSOnumuXbpKvLNMrJ7T3X5HckaR2EupS24
/jgm/Nks7zn8Zzw4yLF3ss7cbMRjI88TJbKVYCzJ3H01VUcmIbC5gAHHwfmc5Ems
dtWELhfx1LJxEuN5ybjuXaOYyEvVYDX1bSpn5BWdMwcw0ESuSqZ6H/pWGgcS7VwI
mHUKFNHbo5FzEaagx2u60k16ujRkoARZGB+akA2l5eRxABC4I4AEnA/vR4uqo+JY
3Eqsj4obKO9CkMf49bpspzVJpCd/VRIkDt9dJ3ji92LLjin3POXFAQ93BwG1VHkh
hh1TAdFNJSs3cWSaNhm/aCuA18ctIQCkeFY5H2IrZyS9zQDMrob4bLXu0mHJBx+N
xMB4n6v/Sm9huVtXHfurIsHw8brUT864qG8VJDFxdVOo95ls0A7JQcpJsnMzbYwH
s8JXnqLYfagV5l8vBO3koT4vrdmnfXAaOI/QZL1ZbIWD09bYz/1IfV5/BFAjeoPp
3S0s5XEgpiwFkf5cFOFP9cCnoBXtUWqDw760XxZORcKWksM5gTr21sHcJo5VHS44
mD9Qwx19w/AYRfI4E0mXQ4oj5SX1iZJZfnyvNRMkrInF4XZucZ+B7Ncf7s4kn9Tp
Ahy67a8DycYKR0gi2LnO/gcNGXN1PgiJ+ZxOuz9wmVw8VJZEDv7Nipo61PNVzP8F
xp/hhnn0raO3ItNJgGdcmTEb/JDQgtmmmLUf72cTIAx9WfnS4R4kWgOd0s8SdQvC
721YVqsE8ZeDKMoa8RwYahLzkESAZfdj7tMZn7WgdYwttmxmSZlr8Q7EfarxEELv
zb3FDIuEqyRnhrWZeIkICn3fhc0mPfHkInr+DjvjBWmwJA1sWTkyaRJWpRXsP7aG
Y7BkX5E4f7kgqoF+3erp44RoFeBWT1xrc8pHUoB/EpJHVUWwiFOWDEvXxjgJ00sY
bo8LcXseBoosHdWLLe02HaFg9pxd1jCK3u79LczQUhWhZQSPoDrhOGxIZHLMyyns
dsJLR6Bqu0r9ODjoDh1+7Qwj/QPJD/WcoTqsUy7ctiq7ofEsOBLFL5vLsdyVve0c
ESf2D9J+/QX2tp9KHQPB97MI9Xkdpnpr0zkEUjpV7o16X7RDIzHmerSOrTiNyFc5
HxKrFsWN4JCOopaiMFu62cyJv8zFnHfnaeTxCx14mxYS18SdqC2zJEQ5Ews3xwVI
3QhvusD1fIbDp3gPLDOG0TcR5ZcKl0E4aRZo+nURY9omo7wqF/WgzmgFjYRf4MkJ
So124K8hP/1sp1bGouW6rBrl07s7evZSF8XQZwaCmm7nSJy8uP3vLkC1w9jq4guW
JYRFw1TtTlfEuQiwufilfxZqQ+KICOiw7gcOJj1HNB9hP2PLFQIxcavhtA+S5BcH
GvHOC451YOvPCbrLA5HWtviEDD+CYv3h50CxC5fEbsOH14Y8SI3yQm/gnL3SwBe4
fL4Nx0hMktO4hRB1l0plqwAWJNAPJ3M37OeK2elDjSkFtE2QujkeDFH5I9watKmc
tyOoW/x/9bwdPtWlIf3zODT1sfNvUvUIsCFveflS+07vtNzkH/fEhQWkTulZvEl7
ZkjrUYBRod9qPRG7+6bxD6pVbZ2mGlxdYUcZwoiyaj8oL6R7yKWkOJdPCEObkxm8
qW+H19hzxU6iIYTV5hNvYMwI/bdHYuoZ4x7M9/6onBGoWp4omquvhhOuPcXNmn2s
Oi6NstGZ8NDs+TRcgR0CVzm9Sy03mnalnUk90jxchJL3agKvmjF0Tu2X/+e+JrGv
2NSnto7TT/gFCtm9Esni7jJFIvXq45Z64f19zAQkl+acf0EpEBn+Al/OHghoErHP
vVDJBEyZDS3NbujJY5idibJNJTfsmgNbQXHdhtzZOnxjkvt1BprIBKe7444A3HEf
jwMNirKpk1SZhA7WBVc+Uhl/4zJwbIMJqyqN3XXEmS6tL5eYZo26ziMKs45kqG/C
uWpPXOY87ikHYuhW/MNNRaLxy9yXwSl4buEzQjz7bmgKnL3+bmOSd9u54zC/MzQ1
ejYlCyAsdNS8I2516EmE8dKSKOJ+i8DZZj8W3t7AUzQRlzrHAnG1vSPKvSCHdqC4
hBcbGk/HWXb7SnV9IafJPE5aFa0XgGZCXDI0E3MRUHNtuiYiSX43w3VCkpvU1HXS
mqtf4Qst8JMjh8BiQrnK0+3NwLHA8z8ewSv3gTNlV7nh8ZLUkaSk8QE0m8wCqrpn
pExmTiUM2Vz5RByuR24TfDUtYdSOgllHjOHqh0HHFIJ7yT0eeVPw3ssODM5lGgvU
sJPnXIA3un0ZICIFTuIOvpmqQLhIF8Zph8PUy3JVIyuY6ThHBQfJJud35jEDcwL3
LTk/ZMSvGLDac4jN0jcormTJQ4NqWzsF3yS7Myr+keg5lmamvc61fU7yJil6loRc
aNxQuisU6D3jgEQg700FMNwxqK9kvnv4HK37Uw/DSjTaC1jg1R/gDGM5zTOA8aZR
W3DAevRDGVhgkt85K9Z8nxWOl2YI/DGZt8j7Fu5YzGJSATgOiz3nowbzt71vUL1u
f85eFuecjHDS0iOLVjhdL35FbsVFHDaeUVkhFdAaFguCwWkKrWhN3Qah+XO0bW0P
2+w36NmTcBtXXTHUbb1fe/CZMUfOcpX2BGXNR/LjRSCBPnJUkEGXhTNObQvGlwXD
mUvC05s3gHzjqXcwJo6euUcJADxEnXIIdmFHEd3GB+g6xkiLdsdmskPq28V8Azpg
xAH//0d8fnbVAE9RiaGVtoXkhYwjx70zy81plSVXXbEMlaT5Rly3TwTDq09ZUbFB
mUJs3dinwlZSsLr/4UgrXIB2WgNp8ePB5/xz1xRIMkTkFwh7U5G2w8AwXqf2buHk
yhwzXB2LdxR/HlSTlHPNXVjk2Xw3cY743LnDIxVLrrBCJeLUSe9VyC43zrYvyENh
Y5zfBeBC35JSBrboEUg886H3znQEU39nL5lOFAqCmnWb6vIdYooSUp/2llYOXCdw
zqH310DVkLGSNQjQQfkXs2xfwxYbvbmQgS3OvHX83+0e+hwM/FcgWs84YhfTIkmH
xTaOEhK7Wh1W2SSU6YT7aUxsej2OAQVJTZzgBqW0/Dsy+WJdJ6tjCWDO45ECDCNv
SB7C/3RHCKynVjGPR90/9080TgKZG602IM/o+la1YZaHnfOjizjIhJriBv7S4MCv
ZEUCfXIFjI7gU8kubZZv4xEXHFSeBjWNtcHEsfaGC10Pvej3R3p/PdIg8G/wwzj/
FCMLojMIG4jlVjfL3zfWlLDCGZ0cMFqKVNBFwUF2KAYGswRzvGpqH2+j9m4+JjoK
9IibkOr5wm41waI1cvKFwtFJvmQoTLorzwG4lw82CLVzKrKaIHfTcbBcfZ5PfnpW
OP/lY2S22GscPyuhIQXPQ1MF7SeC3EjLjKpuMrsiDs5dAqQYsv1QWvP8TYEccBan
oiX52mAaE5kj31RK1qcYhzIym5plKyZRRKoFP/Wt/L4emyMNntVgmeJR8bV8qL0U
pBFWM8IrH9w6Qgf6UsrFf0TPIUVuKt7vFF4xNCvy/0PfXWO3o3rQuXHqZaIHbIBn
PpoaqtIWOrflm5DM2kk5OvO2vIpEpX6lYEL32c8UiOYIFBHeKrUQ0ejZ+AgFhez0
i3/AhyH3M9rMqgCeRZ0JkKxju0XE2OzOkEcGg4i8SA0InX3Gjw/DfwLVcgGZuAwY
7ma1urFQfw5j/yvIhRryCPTxxrLM7C4ZYvALIuIAntN0KBDvpZO3oXBaPwJ+BWEW
eJCtL5a0ifD1tYAtQAAZPkC9a+lKAV0Acf/h6NOpJPlOUXSxDZO60+prAE6M7RwB
/iW8ioFNHVsdCNRbYQxyCsy96OAuc0nxFTt3cpmJXq8EQxZcokoKBeEsRif5MSni
UF2yXIw0pB2pDxGuOqiy6YN4A7oEbZHT2Mt9gMS1KnnFeUHDon4sKPbV6rbw5gW9
minwDvib4SuUJxBUqiKqnv0rdllRq9RoUFPxUKTS+e3tQ/6pRzow4iBatCqkIogF
wDnZW8+geG5Qp5GQQaniUsN65H3WtY2LSfrZL15BgBsbDfVj16Yj1y+C8xlsZaAL
z25Dt/y2zrAlCz4RGJhNEL9QmLvIHjjYEVcfa1Jftqy/uc14ryFmMnxlUozqsI8X
fgsUlb3dGTc5nn/tC7b1ueqlwTL0tMzLaOWFT8dmfv0XfBGCpQedgBnONOi4jOyo
TydrVP6FCVjFb7OCQQ/ZChd+6nROF8Qu1yl3n7Zy1RDLMBo+JAytD/8+d28KqWXU
UpV/QZTvZctaEqXbNvLcbX7mDQBE4en+r5XfFJ+Ixegsf1k17jaTHnS4FOjkjE7z
Hh7tqYvuQzFTGhvJdAj57FMH/KSDUCMOA+IiG8hXJ790y1dRInuu/RhBxDGk2hZr
GsuzgIanwgTcHVq8+rW/jp/PZfI2ZL+UTHworOtQvVkCJfU2eF+RhU83gB2MEBes
FKfDbkbjiyX65SUYJmgefNcZ8Do2BOSvjkKxvqTKEKKPsFIV/om32F58faOXju6W
1Qbd3wU+opI0uwFsFbfTv5eeDrc61hEa+HZQ1NSeiWMCh28bn+Q5UOb5poj9GbB6
bQEzfve9pJxqgQ3e+nkV8cpaEaOrGSEIoHmg7ywLUwxP6zXJMXRHdiMVlNtiaah8
G4dL9fjiliMnjbvnigDzWh+dBoRPA2mrwjWQOR8Gf2heWHAw/KAYVwqlWwFDscQh
/XuRal/kPUpaeB1bqfjiWBmTJmJif3/1A73a23UXjrwgMHjlsuX4zH5DXIbC1Dh7
1pUQ3W/Gwkv3jUqq7kyyxVGleE/7o+Wy/qhLjIj7DC34AIHZb/F4ynLrhTv6ujDS
EgsPEf4PWb1BJjN6vUh7i3ON/+BILMS5A1CZId2uD41QUjKejFhoBzwl8QOPb9Ny
9/HiOfxwgSXO/woT7SpQAyw0IGKvp588bddFjwxF839UHmwiaFZsPS/sVR5kke5v
KFqhT6v83mfaOh7UkU3N4Fr8SWxi00XkuhNJzP9BNnWVJYLm6CA9bCM+H9Tz4pKt
6ypTAsCJd3954Ly8CXcp5/lmJeTeYXB1cwcKcV3ysw6r9jos2g9C5rg9t/u/j/9u
6oHKVT2ECCLXuLGyXjNH1FXfpnAxzWoTyKu8isc7ZX1ABQGkfWrVcMoe6gDDK+ra
2s7QR4kqCQu9WyRvrr0SgLSIi+oT8KqJT/ykYkoL6FDFrdEza2oxj6W82ZI/gDbx
6EmTQwOkd8D7f4PlDoZmFWMq+gylhemWS7CKNO1g2fFM1t3ankR6fQWKWFtpL6PI
pmgbv/VpdWzBTLt4Zz4xLZfH4Jxyn2zT+H4Yj8vOjduScMT6JgpV/yPFbhOVxG36
U54AOoUY5NevwVuQV95iCatOkiZP++9MadgNN+SRKt1e9PFrozFdCR3qDcLHE4O3
9by2tfoCahtcsxlzx86XK8yb+vEkVxNQg8NNBl6BCeJsIhFCHzoAMky/3LET+J1T
88ikEpwUsEpXslhqf5Hl2qFkYKadWFk2ZrHolxdLp7fJpAnrpGA9M07CuLaEW8iC
rdxvc7vqXfB9fB/vftlrd73SAl0P6pbNhi9E9BI9C3LLJ09FdRkSB7FZm2oNmsDJ
pLIRmhOLgLmifFJWlkQ7q4Fzfu5mm/3FMDGecOk9eT3xbCR5p+71OmgvCupjA2DW
Kih7AzBF8rtYTBO2lb+tXUJQqaP3zldYbZ836bIjBgbZhyFB1XAGa2VIk8xJMPqi
lRwO64qD+7z8JZVx+PnyzWsUG/W+7W8308y3fxNynyerGXws/+1xZzW3XKmr6KMr
h07vKaByEZ3TMzY1lujvxDIHl7R92YRM0e53rebG5GhHWEslpEzKS3JnMKbc4k9Z
hur3jvEWtMhlausRr3bnSVfday6eJuGHth/DY091S8CUi6Qcr8+Dx0WT2WkRZ9y9
algI++t0grDWV+IVC/H3lsztapjnImg+O1aaWZoccA8AG9TnY1LZrRMwjCHIooGI
l98SK2vL6Xf8Dg9MyZTM7NKynoozczodZp78TYf28cnrW+5MN+hNI7C+/+IEvo9b
qFDp+U6FkLx3u/+W9nCqQALFl765gEEzfNqkcgHbhokxgdiklkI3zbNK1L6zvw4v
UC66FgmESrpNr27tbZML/d5lcq/t7gaqy0/9MnL+wsG/AJ1jda3x/rYt2+H4mIN3
ffj9DeMobwAp8pWIT/9xYcb38N54lh3Ls0W23RSE0pz6d+kMVD89BKGWi8QRaF8z
7Y+mjXxh9pbmYrUaCA4ClpXSc8OMrbs6M6LARErJ2qxdno4dVAbXudNLuzgjXzPH
bYF1PhpXCZeBM8MQ4nVrR5lh2WbAUWSw7yV5GUJK37isJD5ir9dvKvUjBiYxq54y
nqrmyC1vut43NLvg7gawmKj66uuKbmnsxu65/iiNvWgCo55yAqfeeu2TArAU1WD/
apQAf1FYB9Xoohmm9eO4S1bgoJhHcOaxVgxliJZ+UwldVgGY5/FhZ1js7g53R/t5
d0mgeA+1P7jVIJjGTX2n5MJUei8gDKknz8Qva9mXITcLS9XsrUrwgr73SnBPyQn2
+YA4gpBtVgFx5YY3hRklNBV8bpajVCjFta7/6/DsLcIHgebEX91lr/CjskJMae+4
0Cvpj126NPS8EFrYy5ItIqBlWPZWkgw96K5djeQ0GL4NEZhzorjenz+jREMZkkP3
XQCTAOhS8VhY/BmdDuEzOphf/7C8Ar5hBP1TIKZYDPiC/8iNjyl1YB83K5MHZk15
F6yz/qXDHXhQ673ve6+JziKyHx/nsckHnCroymMNN+lBlssJpc3wDszPmV6jLMrd
IPjJg9aHOGZS16AR9gQlJin9gyDrIF4w3E/RYrrmecZo3Oqgf1M6PpfJDef5BCVu
0zc6bMrxvoeTLauF+e0mjmm3Iay/dQ0OBhRuw5MYut2vJn+FOoZAxsS0PfSZbRDj
NQse18olYxn7q+qN3BZnZdgiWLzSuFSGDa3UohhN35bVFtub71qY+bk5rSYDvg0W
fxbQUcjwpbo/siFx+xWmfjsbvFxyKXmb5fSKhCVHDY3zGU4Jx+WA4JNf6VZe3nT/
/08j1WoK4tir60P/w0Ooqr4AoPScwPVm+9J7wJxJyJM+Sk1LClqsmyBlMycZ54Wx
TqtyQNO9S7fy32EzVYCdaDD2cFN3ZSnvv2H7SetJYebjfHFjCbIqJfv/3xmGC84V
CK15VqPjeRuCPfSo7Ru0Sqg2dfAr++b0a/iVZJWCDhENNEZGP8LymRKpqe9OFfYR
TT2dFGX61cbuhGZr639vq7CcU11DuCbHpAmr2pi/ALgzQ6fSJlQFp1e4+05Bk9ly
X6U0MrfE2HvMViGDPWaMufdvmNwiL57MVwrFgyN99tSmTWKTQ7SQH/ROVLcD8taC
ekiOQ0tn3bSjKaanldJfp1dEaGZsjYzGwjad+sfsKYOsZ/HirLbBMbaoI3NEWkA+
FPEfqzNdRzhGqbSvrqvbXsnXwzcfYebbrmwVKwRBCFZhR1mzc8Oh3sohPyDnxwjJ
RpSuwVQC9hlcXGzo0CN8QiFdTo1shePfVfZ+ll2r2CwsBZGbLs2Q0gnUomv32axe
faNV2HZZLFxa2vfsua2SuhuN2IG8bBjBnPIcsRUsXcwdk598cbXQhHSXe8V7tNni
LOkkO7vAZ+uSOxTv+Xt8CX2hmD2k+DxSi2LyGXfagkKRh+Z9oH9NP3hmJ68/Qw5j
r1OlXgRCvAoKNMbOVWnVQZ0a+hfUXP7VhebgaWweKtiZV27vMf9t1GDsJQN+LK39
z5AewvOC3CE3q7LrsroszBsMVxfhmIwdwBzEjb248fT5zhl2GD4t3cIun+ZKOHip
MLzavXq9ED9ZXTTWc1gbyO5i/dLQD35UYDXSJmFpvrqWOTbt3sJOEMOIrHowGVSi
Z8FKZsZCFgiIHP31G9UCnNS0mhDwdjaRFjSCaL525SkUZH75yO9UXQKBu7BTEvHD
vG46lChChTN0iFhkkx/ef/TguRHRhGXT6J1ChMrnSgtOTS/B7cYsHM46m0gj75sS
7IoVS6dac519ezKMkPtNTQ75SmgUblDKI7rln83HLx654La9ArWZnk5KFKxKYW3d
Zb2hJktWv1IBl8qJgUOleaInRnLoWYHuQHu95nlmAG3oJx7YoV9Gbdy0c1TvJv/R
K2BVs1Qeel2nFjH+jqKiHv16BeKfmL3wIVmFKAS/FBdjchz2M5LH93GVxb/UrtV/
TEPXIixrc6Dkuy/WxcgtIqyEy0uH75PnJ27XeGd8cWTiu1z3j0YULb1B5Y9bHi/U
UqEzA/GvK9iUf+3y7W9j3hcSdClX5ZhudFkbwKgbwDMxGIWewfl0bf3NrmG2FhV0
KQcSeSi7/Bv1PPltYtG3ieAbM8OIb8YOwUIbI/WpTV4x96BtINQaKtBBKWU+loQK
Vfi0tP8Py8tVy/tujmmOGzJqryhTh5pLlHeTx8bf65AvJVFhIlim7E06/ERuxC06
E9bQdgm6N7wCc5oxiSS24iBRenY2FSiQGdJWaS9JXCNnzvASBSr4rdscpEuOtqYt
4yYM57V+zhVtKC2ItZrqVaK/2kh89J8BmjybSDatJOOtrut22mKwkoyH9O2MwoAN
rapv2Ve+9XxkRq9D1u8W5Q==
`pragma protect end_protected
