// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:51:50 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jCPpwDUFx4ofvndk/aBL+K0tu4u+OCftRFnsOjR5e51qDI0RRiD9Gz5PG/dx0HG2
31pZ3UWmLb4d9GWEZwgt7Bk2liwZdEbPkDdEY39U8/qL6pdvloNrqMMwnmWzGo7F
joa2C/NB3ZSPor61aeP7Lx424EVTxARzhqhjlrLxh1c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5856)
zIfLXM2g6x+iVUbhNgf9L92LqUYz0K0IRlRAobatTLLCszXhPaHBixYy7hbB93WF
jq4H1tyQni7RLAfE/Xg6hLiOkXAlBvCa58PPvljTHRZTr6BPxiv3IzH2K1vOXr5u
93edydnQpC7pctvV57yni2bLW2MTmybS/anBH6aesGbIoYN2w9o+dL77MMf3VrgF
4InZs0puhoX4g/uZqxJAOivggAP5zCLqWlO0tRpnZhyRWTPA6uAanoWN5WokHSi0
VTfagQcFNRiyT1PfFES0OFJCCCKFUyNxO4M6AkLa+13EBnw9cdTANqX0Jt71V6sz
9FGtG7gXC/hdnlUyTM6s5q5p3JDjq2aneQKFof6Pzb6H0gI0OJ18313NLmN8rn12
zdTMBA1X1YIqT3I8+Lh/M8YzUa3mATqX3LojtgTTv0tLl+uHDjftGOjyRiWGNyuZ
FGrHpMJvf3zd0gBY6CUeLwuGXRy7ARQxSufIdgJKl2xd9JkR5Ri85rdvPyA2IA4x
8x7Jv9NELUhtYPK4c/pH19Q43IjV1rUk0e7SJDv4BM8L5rsyH6ffYS+HAyzRtSuI
SYOmRfoPSpMa01XFpxOimo1MkfEDahlydi7llC+YDnNXRSG6FYqXs1V7zAQnpLPl
cDMjyrNu+bPmYe3k7v4x2AwyiCy4GONjjwvNE19DRZQeexH8AsRncx/ztxkhap/V
0T6vGbMyPni6jYq/8DPQCQJlLffAH8LlJlbqgrDrX7DnUftWJ3QAmyuNeykuWVrV
2+crlcYFpuY+E+VlACHrbHUwhVCP4lbxPwlD4Xg87cVpHArvsX+5n22ZOquBQhnu
9eD9pbIYixG5CheothuGUPS4llWQTG6YAbjify9XINJ2JX7VIG03N9fZUbdpKLb3
mrpr1kQiqhIvhxImUBdzCzNlviFflY34DvhfPHZsyOy27vmHG6mkxCX1QTPZ6Ylp
iKMkqR84LicZj7hipNFXAh26LNnY+ixjLlKwUmy8gnOpjHNb7yoZ+gmQv9bctaw3
X9eC8itbnault9zmBAYJJsX2/6pyehxqiO88F7GL4u46P3e2ZkGgblETbs30Exv4
bacD6vVM/ZLqRsqgFawnfC60ZBTrzOl80Nkv8QUZrvGpc9/1ZrAWr570Mxr8znKw
F1l3d7BXb1ul6mtXhQSzUXelME7WlfIFT50gs1auD1gi/Lvk8g9oVl/uDspdxC88
be2OShMOJD8WD9hfaS31Tt//OWhJpAufDG8wBTKop/8HxI6QIt8Z/mz7xsckeK3h
qmR0HhVkEyBX0mWVcdm0ki4hQhq9Jx393ighYfAYn53X+9NMqgatZwxY+IoOU9q9
8J3Mwd+sIiHjjAlbDjrRJ2VO/VC/+ilsrYZVFf9kIbBgWC3Rgow1KbaTJ7Fq2K0A
pDR1mpDQFixeOLKqIdDZ7B3c4tWeKzrAUAfDwxddoh4k2OFv/6x3yIPPm8pBZe6F
ad5bN6TtO/IuBZhDs0sS/oTq6E7T4zfr6+/bXmNepI2rG5aNFBIh+bYRSr+hL/Ji
Gz4wCSAG/k0KgpqK75X5SCiH0DWd7/tIAuUMYCDfITgX2+HwX4QHvXfrMta+ceIR
ezMFPG2guaJPovIkCeTFbyV3FNy+sJwA8sVRb4xCcfi3+35Ol3mvOuF1CmgyFm2p
KidFdhpAJP4U37Ml+6ReCaM0k83ijEuSdCVsip8n1siQ4zfFn7VzoyW+n11FO3zy
ZQr0Ascd5Cy8u8rbPxQYqtwVycn+VC1+AJK0p+PMz3iIhOns3os1EDMlzQshlxfb
cjceQv0oSQAyadWXHIm1iDXsIkFrWXM+hpF2bnkl3Oo9s2tYmxOApVaITlOj8O+6
RQ4/zx2avoSUfv60jGDTBXJgVuw0l8aulqn/MYawoVityG5DE6rv/nain8ebQGma
7FK25+nKrDWQ+nwgBtd0LsDtrUjTz0ErVaHFaYerxd2t5pvF4fbMxTCMUAWrZuvy
4X3z2I3RGfzcmZKaRONQcOdpJ0seM7MzLJK/iqo2tXbd+RxKRtN0PcxvPfXY0oJl
qGybTwbZoaJdzn2K27wuIy/1gzixsbE8wt9P5/33eNdqUJLJrUbKDld243ae3MN7
To5lMoEVq2wz+H9f9tWUDNY505vnevGQoTfo7gIDmOUkCJZv0/y6tTNx/18XhF4S
EzmmDFim6Z3ozCwqy1xvcGemfzyySZOr/YOgv4e3+oaiwjkj414/aWNEDQmzxmRU
3Fohgv4Arf21yuAlWYhamNV2vZtdbbc87eHAxj5w3DmlUEhRk24s9qu9xw/lIKgY
1yDLuh+Q8LpcB2oCs+7oDE8yYL935rOZ/HBA8lp0qYXKhqBsTu7FRtDkOHYcT+jU
r9uu4qVQkivBYi7vUsE0HUR2XrPHK/MoOkeLR8PP6NQznGAXEfS3Bb9/UQwhXVG3
+5gCEvfFpwyIGIQA0DnWf0xhSOapfCRQI4yuA5+njr3NaeGxPwb2tcORo4V1jLlF
80VE8veRsWp1EL0/2vbB5Dv0KvZGTucGw3LxAoaBx2btX9gfFcC65X6VPAvhlV1s
9C3PYQzBdzpfKc5jk8BfbY0yDL2ai/c1Sn89040tEbKCREINUGI1YgCLAfIob0eg
NSnJm05qSp+S7Yb+GzjolJbMcG72dW4CLPc6EQhgPI9hLpaQUqfzYbGZKTXpDcsP
cPSSu90aTr1hvJJo/2GS/iEoWQqmzlwVduHsupzobLwQ0FWWhdNCeoZItAe1oDyo
tBQEft2x11KIp2n2CMpz77LPYjOsngOvw3gkeeZjLfjrzzI1wkTCkTAKy6lYMrYr
gGGzkgnPjOCD6i4yV/uZQKM4/HD90V5OVMvLUGJ/q/Qk1azvSvRZhr3J+ke2M+XR
hvp6p1FFN/BNbMs6Dsr2XHi4uFt6zZ83npXysd5r9Bg8WK/tQM0fzwJ2qzsD9hPw
5tGv3FWm06rsUiYXZINgRzyfI6lzYyoPogAPnq4sZ21/efNykiryYA6wk17Xqmhc
VfOPeGRguNRKQB/sPY8uXz6C8qJcdbnHWSWVk4I755kxIFb+pea6Fuc/yVX7LN0I
fWaBU/Z5h0G29lnJ2iBZb++JXKSRZkajy1lzzQKwl45mXB8PmaaNT7MdAnwvRfkG
Lx1uEJHxtrBiJIkyb/7Q+8AFbTBXes5Pqf/mtd0Djrn9JD2I0OSNK5S3rvUl/o7x
6hdq+Jsb4VbQ6TvVx7EMhxLtetdhfs6FrvACIs+XSPaTD4eWDasnJq7dmEpW5shy
+Kcy+Y89gWDkb/KknqAn6RD2GUTSmmOJft3B2d9h8BeofnCQbmzoP1ssQKVgH9hn
al8TqxVFg9+6KdSDsfJZOsguGBxYDyzeRR+kXRav2dqPqnn/ckzacMFogEjsDb99
DkwWL9vo2uyQqoUFSSI4pSc+lGMfHhgO7DIvfhR4+OSWEHEDntjgVt+KmQjkCsIN
CpTrgA/qbNE7Yv+9vHDG8haoHCxyBLMdETtDk/qcPgiuucl7KraH+pBhi0wpg7rE
V7nBQJMf7aty1+02rEKeRwZlELVFFHhheIAjYFTYInF8TkOUqNlQk7XEf8dy3ObK
sa4qtypYMzzxSQ030oToR/JrquTfb+U+KaRSwlk1Hi6X8o71GbNKk7sF1ttinNYj
9TAsG7gm2TQnzBEJLV2M0A/kLH15uoR9axT+BCmKmlD/8CBlI+Ywp9mwohnw+ed1
hVFs8+YQ86jqEax7ZSQkCpoMUWQBjD63wGqrD+l37R5MeOgeVMUVJz+Ge6yOS8HH
zXhHO81FLvZI6r6C0k83A4DjIPhtRKc+Cz1xINIeamG4SiCJSTSDl8v1FPskxt/H
1n7ioPROKoFb96+gi90hWx1OWfnP+eTyPMznyeTT3UEXhEftfWk3wl/GVuD82d/A
z5JBaYORuGHnSB9DivgaA8rmiB/K509GsolX/CKqmzz8LmKGfGeExdGED0Ab7W4N
bHJkYTnNlvONF8nzPiqmj2zP9IdUUfKs5l3rlZdWSP7qzTvtaHZSDMs/ygEvGTJF
ZtLWdWxCT8SWWQz0XP9YOI3eurqiC4SfQ8kHH0tpvU8m/2Fen+ShtLk8fkt+ge06
YWLFKpXEJEVmls44mOCfSxJ45LMt26g3AoKhmbJk0fyRvlzf/rvZFUxYnFDHogMa
k9VbqCo+bmbvhUO5jp8befVw5vfujXAFIykWk5YWkatb1UnFmqn7kn6qoIGV5PPt
eTyTAZSJTGmPfYkFFkRTbZ1IQ7dmRRJIwQm3MAPHYDRQDJ9L5HbA8u2EZq6//XjQ
/eAwMplUmOrBWIG3IT4qaBGRrfL4mnM3NeqB2qwSWfJRRvFxEaCKBux59hguocZW
hzTge6ZM3GIrFe2ebPAhBRToe7seobtjkFNGLwiaiOp50XHzJswuK82ANYs1KZSN
fG4zBCzlPRbhNHd4omjR0emx5MMdthFEYRu2rfMNCC7XfBjc4wfJ498AK1UGLPVr
AqRuIDMAH7zkLT2NhkLvP8nfmQumUg8uzUwj4PDBWvt9LkICjyLsUnn3nQBB/rbd
swCgN7dikBhKNUM/+dTUhQ5zx316hLX8CMCIHdXuDxFqN9Z9/HkTUR5IICtpf0Mo
74mZ7f0aGfH8Aw21b9S882t0vuLgSZmttqY3ntbF0g/+dhHHJT/DyaKD4owuNKa1
TNtgKXrDm0ZaZlzjfJTRDQNkWQHB1wEtiL/9lsJOoO10vteJ00HWEhBWrorKqMXp
w8o7+8lInReqF40uAblb/II+ifWxUnd/B/Aiga/ZE+FRaeT5mSWjANKqF3X1ahWb
Y+/c3lKpNis+FDHz2NZMulgFVHDQXdkv+bvHT5aVp3MqqNB6vc596iPdyZrM9NCu
zEys/flCM3fi40Re/d1HViakH+N1Nlt0XNsk5hlRSLsju1AtNhhHLI0a16RNjrv5
zOFUSfO8njDtZVVMkDFAHQGE+vXirqutRiBwCXlukujDXQdOBWV0EAu1m9VEcawY
ukBgG/z4kvuFO/x9jxS0P7D9iQhZc7L0covr5VtyyzQOGj8d8UJFaZMlNRG8sCG8
vme9qA4R9A/EzuX99F50fJR85SzX57sEUPHpY/jkc0UeZOXAut7ApLNLgDgNAO+N
vbyRve2by07cQzfO4VEP1v5AaNpK/scnfNGBHkLBvcCps/WIirFfjNQEUNsyysmu
aNFgqwEcCXJwiNdJpRpcqEVZEgRDMtqbWIxI5Xi7UJHJcw8o68G1Rf2ki+ghUF7k
tE8EZGeJUbm8qvhicclhC019Q7WDD/cioPb9qvfjSyiStG7M9J/t3ZbQ3ZGzDrAe
ZrRMOXM/nyi/JzqynSvjNaUNoBaRWwQLdxuZnEIVDHdkLtvYWcZ50NET/yakm7HY
4T5f8yl+GY2jzc7Yrh75JuoefrODtYr/aazKbDH1/WENXXBza7rSZ2MmV8QYiAn2
UYSijT723qiRFigD9lMsHtonaHXLYrRkKNnNeQCg0zLZ0kDi6fJ/5fP/YhEpXFjA
t7rZ66mHCN+qyV0TZezFLnjPSa2yVUuv96UtHqOUGcgxH5K7hObcOW6T3lWHvoMt
NuOjg/Ih0SAE3n5VFDWtXlCOPeif2TU6B64JseVUAt+zKDyMwLLjJAIcELWPEAzW
Pi0TNqIUab3njIm216iq9+uW41KnyeAf2q5EuQkRxXYvXYJmCWNSSGBkfx/TWE4B
pqCXXSfbKYNGiOgVM5FztylA43DzWuuasG09PCGpTrpOFZZf1flVaett8RrIEo4H
5Z5TiVamTe2OiUoi38lX+vTk0orsmj6ppYnq59FnDnYGVNFIGuJBhwUKUENtaIa7
JJ4pRgpvlOpNZXts0r/iNekyV03pKYOgGmQ3QdMsx5B741ah9wjE05H5j/rtglM5
7raOj4WARH1zDE/4Z9gbnf1o+DzAQdR8ypieujmiZ6Npnv64PnuAeS0E5WkVTUj8
rjID7XR5NXEGTEYQLQ70jOM4ddWLvqSgJlUnNS72jM427sSiwH4WjN1/m8/A4kT4
kYXCj5DgTxeCvmw0kni0z+PoFsHjQJxXfu0VEaf1BAvc5ciJio2ShtK06vnFU1Nf
iVNeQEo6MtCft4MvQrMzE8cUh8tQtcKMQSMJ91JgJxdzP1BmiVrlgK9dwTqa5rqk
htz9kk/FcIQYQOYG11HJQVZ42gcZiVzA2SWgAtG4rgdZ17puERHbqE057sLnGhN6
Z/5KaXBVjzshgqcXhjaAdyip+VdtqX+Iv0KVJWvwe/RFoNKK2g20u2L6BBa1hYwE
P+tFSpCjdIu+3/ESILWl0FLVexWO8BypTQgxYnRt6BVWi4ZS5WSzb51PDIp5W7zH
N++eixL+eLYC/t6vwPZ7wnN9vp8Chu1QMB7bcNBfb1GcRK6kBpeO4uucuJCoLImn
Ix7LTgtpVN1YFRXVbBWVF6S5r03O0p24g2lnnSr0O5T1l3NTJ9Qhj5uGAtQbzbdc
gx72wmLIo4oA4+97ZqkheVUHXkDyjExtfREg0Vq/DKdW8KaXVfNx3bo8tDNWfUPX
SodPNmCi01bISaTjEdRjjXzcqMsvOE4OrU1yybm13s4Pq7WyLLKxak8oQtOSPr1J
HD3L/k8s8O1J32AEYGAgyxzOgD4XjWJpIbz4aLkhdW9iclBpP3iC9NcYmmzlVayB
y7WmQ5LCTZCzOv84w06vecYYQ3W97Y5A6ZXeryR3+cDY5Ejy/H6rpOJjq7voe+RE
IcOO0t2XI1IneHeuAWdReyVjG05AfOh3ezInT4kqTk7QBcTyar9+046fxQX6bxug
4gT1cinnhegXGiW3k85yJ9zuwHrIDrWsdIQaRtLZ0Olj6bzgQHAe2TM+DUpREL/o
OJwo8ZcPDrsKCshUcxs1C4PSsvpJfblRjwhzV6XFZPX36dlX+eWh+Zh8HqLCEmrq
B+GkA+THICT1P7sQE/m3stp1BJkOIZOwyfuWmBthB4p71TxN0n+o5jIl1Cq9ylM5
ANVCm8tEstQW39V3qnbd8biPpbK3rWElpv9fOG9fMUPBwEbbAReQ4j7aR5/3t2bO
s9R6k9PvpYqvAHlHJF/kvJGXLUgMcDzqPZ2Kzf/z65lCyiFXqqC/5rj5MdpdQE7z
VqLIFnJDbbbTGk6SghjCyqNc59dSvK94QdpdEhhSOD+KmEhKfyetDSR8kZN2XVQm
8G+aLS4w4K1EzucjuSAsGNo3p/ve25O3bOwuRX2Pf0x5QuNC9bxgNQ3/ABMKd7qr
KdSGIH9sm9YOx3PHW8O27htwA2a9HFnKwqARrSoHr9S8i5nAEVAaIOSKSUmW/kcD
kUL4RfAoIReWolvW5r97TEGa/aT8ZUJQMW0PhxX34iICX691PDJNGzt2YWeKrntL
Gq/p1wBaFkrutGrN6ifrCTWMSyz/P5OSlOquwO24cSGc7eJHuhLYfP1O0SYFSETi
eFL1HJdMjOa+dvv1l/3hQNA/5zaA6l++/PRDhK/jdUcR3bPYfuk6vzmX9StrtsAa
7bRe8rXn8Q6BduqmpTcj0OEnS4RIB08d6MZHpy7xUub8kAni99HfvadUaReZboXc
h310PzXtd1ttTCLejoIIy2tJWzuusQ2/YHaSqiU7ziDiXaGUsnfODiOrkmRU+mzj
iUxN8F7+1gYCWr5b/UAhK3qRpytKzSr7hQolqKyL//fgWZKxSeS5zRSupl0zgg4L
znMZieNWgQM/p6h4wY5XfoSQYLu8V5p7fpS+4IPxASHjZIfaXl5HX7Ow5NTjePAB
fOvuUYttaLow9LCyx0J6PySDwMs1bpXpyzhSe3ngrVXGSX1bF3i6mb99YmP48Ip+
`pragma protect end_protected
