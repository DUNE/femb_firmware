// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
fM7uqi9NkhGHNUptCd5hp4bxqBL5ZboXsudP2Lat7T/yREn49S512cwKtStB6AXPqpvhDTfEFLXZ
5CpJtrtbJ9FdlFZeEkHLdOrMnyL4j2iZw0AwiPLukrSma/wgPexsH3F2sg4nIVuSa2ykrXa6CcHU
N7EoiHn7mbcfqZE1mjjxY2e3a7pZN9l+yaulN6JsT1E4vC+RMJR+FIYUx7SiJUHfB7tz3dc/4vfi
Cjy6CIwIeM8n8gNwIcIPqTSRd7VGaHX/2sqCdQ1fi33RfZaIoBqrH6pFu5/YZTTSE33aJTyO7f6d
B+ECaaFV0EczyAgfahvur6013/haaPasdP7B0g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
oT5jknmReI/PkswzUZaDwnZjLA9ojAJzvyOjAynTwFVe4GW/94oYJZEzMKxmYMwPTAHxPzS7VSmU
g9olhxWf79NynIeOEt4XDPF+D7lLOb1JNdla1MQLU8Hc9yy0jnOfihmxZb0FiR+Egn26tOgUX6Yx
817QgYBnwPYsXbmP/hjUA3DKh6LRRNf0BFo5KO7AsX0M5Jc8kBGVdU9bG3X5ZfyQVwaLJqDjVH92
15Xc3JTBdtAvX3zgXl2dSBJ4AEWEbejjfxr4xn0AXi0W8FkUE0ZG0ywhLDE3UUvW4mXPEHEsnikj
7ryD/OZSAX1zr/ia6PGA4uJ4pc4/Gn5ooLArNs0/YAI6XcMNv+rsxwNQS9lxYz/wFB9aydb/rP5X
vytQENL24UeMyIj+37j7QP1mT+naSMWcfNb9f6fd1/kLYyUKNYzTmYedn8z3Iab6s/ryku2D3brK
Aw89ObON0CRcZbKRHBkOcb00nQ3uB5xdzNYABWAaZgyW1lTbWAQXuB1BXoH6ohRwIFQWTSnTocuE
Zs8MXFdblSHxLUv40LvlOxQhE4oWabzlTzwjGJsVIj4vBAV0sGOo/oKoumIQAiC2Iw57eDWGmdqo
RNxx7GWrU2ys2Sr8BntZ0HLBFXIKCNrnuVAKpmCRjK8JE++mGc6HYn6feuZzHUnlguwp5Nj3mJ1E
YGjmo5Y2fpcICsTMv93w9MATJBR/gyW3Dw64n2jnZNfNwa4OzgcYOF0Jq2Q8Zpyr0GzYaDfxH8fN
CtbxtBUIv2WjfESKBTeoFWfEsZ7v8d0WIyrxkB4rJe87H5ltOosqXoaout88IAZPRXssMmj+KjSd
PnaKcH9y6iQtXTjt9gsl61BTsO+Qvw+fYRSAbuUsUxQBMnuWWF8B90lyH3HsGx2HhdtdA2DYPSLM
x2f1ADnXygephGYyNRwCIrLceAYhPxYPC0D+EKRVDeRwZX16n+B34xUdz8uocvt/Y+WDhMW8bi7h
2cQCIY2iTzMY+nfy2tIJNGGCf3Ogs7ZWXVtCSKvBDFzg5iTsm3eHtZSuv+BmLsuZSFHpUY7TPNBO
n2Vh+SpHRDlo6v2IA5XRvXohE9nCCN6iobL2ufUNhfiF2JpxKj8hJ3xTes5LfGqMY5V8ByhIOM8r
fWqiqJvzuPUHkRlfbWzgLKPsTcxI6J86ZkdXZh+BhQRDWSq6Z0i9ZyXhEYaE3ZRc7dvW88i4Grxq
kk6sGAeVaM6kJDM7X76Yi5U7Cevlw1mhTId8tDi7NwAawBJLHEPIcQm3WddeFXqZNwEdV5IU4LuI
rxZe2nnaNDADMAZsXparBOls+PTZsybZAXsK3X4Gkw85rUrRt/3uUFfbG9FIA6CIZHb0+fFDuwTq
+UpbnCQyj1WXJ+9CONlhnIk1DMXVNbM4BjCj1JYDb7YxGU02RoGheW1rRizb9dNXESSRf37Ypf/5
k+A3OjBXqHANwCABY6vSExafO1P+KLoVT91XFSpQ3OKXSzVewi3fVOSjTK3k9yoABjQRmtqe2DRL
ZSobDbLNLbSLD7bsjCVOXjgKx2yTZYcWV7+jTJ5QSackW9hOwg3aJsZDrbX9QC1OzitSyICQjfWJ
JQjwWptcenRe/tLKbNWPZCC+I+p3hL+Ops0nAXa4UYiqljJYwxYuXFspIC/adYPNsYs/3P4zl6xA
WsKvP/vjZy1sGWgccK8NHuPUPK2GWae+8R/rcvHOPieojDm2uSQdVrsCDQpkrq1tcEiZ6ASjV8Y0
/OoMOBQz3NqSW9MDzGtHoHdgpLk/udTPvg0/bNoNCQA47KgbMyPwTuLYykfdZ+AxmECDtZRC1+50
RLDaaNg0VoQfEbamPPaM7i+fFB+lhf1af0yQ8EZcOsQUkTk7QDpek9RE7HeRxaDJwSRVxdnK/jvQ
dcSHSNTEI53eItX80sUB2nq4eePfcLgX5ucbErU//++OuQOjieVpLKu1Bhj6LnueHEi98kJcOR8w
vdFzcByP8WurppdihzRlK/u2+6cRrxOwx0ReHlKP1LfaN/umUKC4Su17tyjRlmmWP4Wj35xRlTxZ
Thzzvh83MWZqnc9Oq36xncL7LwqzUgqMKoMLlGQzVqAXEkJuz5yOasHXqBCUVW1iyIoLdkXEMVrY
YHQY7nZhFfvUnd7jpDnVqQePA4XcfnwtOFoL4XgOAJLu4by1sruFrDX7hxxLj/ilmZuIn5j/v82A
sStOtkH2nvLJf9aC5Ayf9Mmk+RS0ENmTzdZaxfdUEEKBDrKBc16Nj9486vZQhEgnR8x9cM+qpDRc
HAl1WYHZ4DrR0WWO5j+je0jnbAJd9oHWsnz2xIhCIOrJH1IhZRqePs7KIpdeP5u4oFj5rSOGqdBA
fSNQyyPVKtCzu5lbAAFdzUtTl8LcziLtbBvzmsLgArSOYp0OZentYqe7ldzuSjwxQC6yNO2Fgcjc
lUSaTDE/LKPzy4FINST9oIuSXmbmzvEMUl8lIs7cag8wxOVc9DaDkrDjqLA5q2ecsMiRRywLHnaP
KfVtKQH7ghb8eS0yDBbiJdLSx6FZKqBLfX752f8w5SSV6KBsDVJDg/JHy1HasmyrSUPs+IUPobhi
LCMLSuhVrlJl43dm3kvnRVvqImp21aYJPJ8gZKcusl6DnJkOCJ9jTruStX+DzILjHSwaZ4U1dXyl
AVbyV+MS2XrQvFBQIhyRlKNBASDoceWAIPE+dLENBlgydzx222qvp7l6eiQ3PvBKFsPKryDq4eHS
TyYQ/NJu2Jz/eKgaxYR2GW1WYFvedqmka4/9+bBZnVP2sUkeQc5TrCiq9ouTApR0nPGUpiYZRTte
nxP7yVE5IINqfVksWjkr6HFU7ApTTYpAeRXbQIVSx6OfdsCpfFFUWm45Prn47iuAeTL7gs5e9hcJ
ipoGladOnN0ACdUWh/CS3KqPRdxEnhahOI13qkd5RzLfPFBftcRf1DiBc4FGbkA1g7eE/l6y5t3V
W08W+gY5TPnfHz+durE5CEPikO+Zpz1SKDlWGV/LtuKKfA27CzufTHx6/x5AtITPWyhfQ3ppa4WN
SafMmVJPoaphx67c69MD56IjNK7xSVi2PuGTGO81s5u3PCysCExI3GCgI8CCbXRQhBrKphGICudm
8gjMqCEs7jkDwQN1c5FJXIKZzEVOCiL7i6xfWIxW/oZI+qq0JbqSHhpfcMbeQ62kTqiDN22iCQgw
o4pp/wlEdXBH8unSiCmoE1v6srKSIQw5QL7OMsm5zq1lG8hSXzJD3bMOyXka3l66lfr0O/SRyb6w
N8HlsH6wZXz7W9fRZIbqEBgirgTs0XNqC6m5l53P6PXDUYl7XCUo/jdB0BtlBseFMttBKCLcZkBy
m72yTRLwRYB7mjzsLre3VX+kUVROU3fpTXVILWAw2MxkQfB8N/dG83drsc9dMe9gSCeN7RN5Fu5w
fpMf91695sklCpYbecspeooP4zuuNDW6dlNdQeJtYNRCAGtb9sl8uP69wJ9TayLGKmEdAMMXT+Pz
Tew9o1IE3KeGTFg5hEw5rSnlnoCWiA/If/Fetay6dm9Dk4rQOppJe9C4G1rJtJctySmZbqgPp1iM
SBs5M2mg2Mmb4JWbkOzCnyWgTh937pHRFY28aPN72l+BN1C2IJ4jm3Mx+hUK64XaRfZ1cOySxX2N
Y8CQnihHhtv5o/P8Kudwc3O8CipahzVP9lfpM2aWb8C+Ad9E2lp4n4zXdboypaRUKTJw2ZoPS5pF
ZtKOvNYPLQ13t3m1acRy/k7L7m7uuePtsDhHcDXCf/7V4moLDNA5EJtvhcY1s+OLpP6DLGnbooC9
722XzEW94K9D+UxIdh8ilELdUyNnbBL4XgEFCcpHOBkhvwaLk6oeCamD9Wibo/cHgRJ0aXv/YR53
B5sdpTd6u7/YDgMq6/NAymRJAkT1Vimh+F34P3gt9x2FLSyxR+2Ad93bV0q9FTDAPMazRYYOPsn4
WPwnOpfBQsD7sKeLDHo7eJioATz5FWy5tWK0203+fjDIgfJLD4jz0jWEtd6ycpwmdzUrztFhBpNA
KZa+9/eaZh93VJPbXzsrOe4sAaHqJWYv/4vIoXenkjm8NFbq8xV5wsmg5z9XAfZjPxaEgI3+1XFN
HBOqxpg+mMhUm/2SYfWiPtj4+QaPICH5UegGTpbU3y0TOuGpRuWcrTMmWxDcvn+J/dgyqHWbyM3m
EALUyB49tA7eUNUfD4uF+7If6rIYooxJh2JffLObXKuwFZDpKrKgYv+2KfsT538Y/bF41+8QfV3V
Vzn0j4pN9HiKTJB4TxeceIwTVgZjlbvN58Bonu/jJwC8vGEqPQIAc7FeWGXbt30DrBfV2yBV0Xml
cbImzADe5K1CDccA953tauQb8ijL8jeiGp5jDpHGAKvOLOg70J+6luaJJMCJ2Ssuk64nl0cdhZah
2hABdJDUsAOz8KmA3cvO8lvANt7AWLI7816NEcsbfXdDGzihlqNsjZtwC2LWCAknuyYw67g0yZqu
bruwvtF6egSXJ4frzzuu3EapzZolXnSyku3qlw6H5Hcn6Sn2j4Dg/Hcb7uRJnpCN7gqwbqAN8A60
/gcptpmW9vUS3xVCyOcB15SIuHXivXRCQhLo7dShbczEHwubVEZJoCN/7xbAyf7GDnax8wqyGv2o
gNWh2PW0IqIifdMdEQ2qCegGFEyqSahKoJoaulKv1aBYU0+6M3BEX5wIGCIelfBOnOuPcZHn0DIq
R2bcsRdftVDDppoP1WrmnI+pER2ijSZd9l+6VqwuA+ovV1+qiiJie+1T33LTqdrU9GsT8zvSQrb8
DgBZqhCxlSDlzvCM7bK5oCpLiVprtU8mczcO99qDsQZAgAbLITPq6rHjzlrcw59fynrBJ69vWOMF
YixPZNzR7g3wmnGHU1QSDTj3dZRlnN2ccQ90H4x97lEB/F//2pvM/DiqArVk5QGOCo2GcLHe+ECz
cu1BIubtNOYOSnJ1EpMhnKRq/Q1aiXn7wlYfMEfO3FYLAieVPQ1j6lTTpYKoaYAoy7wZYZzbSZC5
7m7BssSJa7vbPlvhwfwigWUIO92whHybHFhRj2UqpzZ6m8e/av6Nga7Imwhq8AoBcmm8ZaOMBCFr
uu0DELgiGEOlkTGOuYDq7XbvLIGNOxba9nN4hnhVZT9uTWkqAcvs92/CDRoumRQ67W6NcmKMhSkA
ZI7jupbZpAu3xZbg1nNoLp6PrJFGw5OfxP5NkS2KFm3xKre4ki9cKUKnOKsEld3hAsmRa41v0JOJ
PVUX0oOUdxq3Ah0HJQD93YC8+JAiVPCc7XqKgBVfTHhvrmCg/U6YOxY1vNSBMDwzjbd/+UHjYkm5
q4Ic+Exr/50e3234/WUGUoW1u/8THeyMwHTWTAioHqRHvmGT6RRadoLCsv8ipvrpM69KVVkPzGb0
SU4/7Z54+RLs8FyIVkquHNYEnidyhzM7nazaJ4xwOxApxDcCmoQsG1ln+d3NRNx4GjoLKjmV2RfH
ttJc94GLiHpx/HeTTWWz1cPkKjqVbaZPZeA7RF14l8NbjgyC38YASqpqw8SRs08A5b7tkOtSKnvt
BHR5vcZkl5BtQf5zCr/Rr0fPeKghIfur+8tNo6xqfx27gyskrD8AUlONs5WeH0mzWnXIv3GtHB4y
/+L5cPA3qupPZttNqc8aLx07UmNeIFRO2ebDkeFYeJ81E7DlQG/K260cSJ4DkmcCNxVUkAId927y
HXgukvMs5gVBQJkuHlj4de1jm7dwhoVbMkyq17uldZ0aRaHHLAKl0ZCXkyVzcorj2UJ4ti47J9T0
cJ1diurDMjj1q1VhHUSLj7ylQ5SdIA10AQaIjbXJ2t/SeQtRtGgpT2xsc8gWgF38hdGcPoizCkFu
KTDzLlFxUOpqNGb8YgtOoUCyLcgRoOW0KkjP2TxnS2BySKKMMH4Sy8qKqCA+Zns7eJf2AOayos90
VsIxxtJHgqm6Jbr1P9L2Mm05U0H1QTD7XBqjQ511liHs3Ks+XlMYlMFJGshzRCgibGGoqrX+M3z5
ts8KtbdtzxjVu+BhXzXqi2o4uzDVwzTkF9lG0kmnhvmQCbSYQxMuHdsMEPBUzVz+uJTmFxYeRGDv
D0VERmjHER1K+ya4zyhUNw2RQwmo3gKA3skv7uEUF7SWmDnvWWiaOU8y4oQNc/gNzPkbBxNB1bOB
dtdaBHjrcQswtDEb/STv7GA4JolTosmKXlU8wtx4TWuZddV1toM9SKwkqWojjlcGCk7744uaCEHn
14eWP55JijF03831cInuXTWp/f4S/Ls1ncHQZ9su7BhkXhCln3JrFKSyaYe0Wy/AIWf+XS4W8WZU
ZS9bnF9z47WHVnmATOdGTobnnZPguZoDgWVnBRBuf6IAoqZydjDTeiVBHrowTlq6GzRlbOBNn6H5
Vh2w2FmwRAaTJWmZ9HC+cB7svZAJW9xxfWwZyiPPSNa2lDPsEfC+RGpdeKRrcdFJ84I4Nd3eqRO8
MOgEXqBxQA617qtgpCHkv3MNi8OzbE61QbnM/d742eKQe0mS82OrLskcBAwWdWgQDQIajL2Cb9Sm
A0dWLxKxU4+Zd/7c30bYIcv6EhdMccnaeXkq8rmI3qQ6G/sFesTNJUw92x2koPP7FomwinFDFD1W
KFcAbDkfYIosB4TrfeLCw1ylxcu04lfIk/3Q43bJvuiGy8tBUDOeG+o3YdFLjJaa/cEa91O8kEUy
HyLC+g6hK2d4CrMYMAZ9jitV3CyVrYa2KX9HlHv9OBM1p9lhT650mHHgaZtMCHwRticVUO6sj1Hg
OldnPyoAalQdAJfshG5bf1yqDCSLoQI2De43rgUGogGTJ9eBXWxvxH59XyjWRQJaUfvEMhhb1m6m
pA0bEtyto9KpkREmAPFbWOyWsT/HdpLpKWdK5VyQtVsLWFsEMMptfjUF8m2yLLckOJrkwltMxoWG
ivBJffjRiLiCtmVUbCetYLHC/wFoJCIPVpwxaXw8doTmMxQADWSbCkLtq8tGK8MABbUq+ZByWZUn
gbDGJtArHKh4b2JThXAA5K4r5TqEsgBzBBjmJVQ471Pq7GdqI2s8AIJZt393JRuJoXw5sfW7+DCl
59pD0LF6zG06VjwpSawowUfPOwRsdLHlkUK819zWKaVeWkN84Ps/GJYwGsJlpeS2S/4Aualou23w
7FKTYepG/SOMz8TwXuv/w5+hpCeID4YFZi7NhhYI33rBrmjUp46wdipuzUTsOen7CQNo0YQVgbAU
yIcy3baH7szAJIvFaxBTIrX08XB1k0pJeyEIyQpARgKIw9e7Q0Kpn+3+yH5RJhOfdPTfPCn9Rqk8
1MvkqbpTQAD8+wxvwhrCp4P67WkvifLZAHCaf6I0e5/N7sa9bu5spdD72o5kTB+OxHmW5YIM6lKU
CUPp9qtHzSSEUcaRAypkNYXgDavrpvrfBrEPips+SVsZYUI/3RFlzntKigVxZR4WZJopArb6wQzb
3+KyN1jtlKWc9KS8jiyRPOtN2j0VgAuqocTKqUvvZXRXO1W2WmChgIB2lmDVRqecwCR493g8hoFm
AmxMi/O171duPMt6hZrvGqdNKlbj62tQ59wVfHnQNQUKGb1k6e3uaXyjR2ZJDn2B12+Mpk3s3Y8q
xjKYskjVzajsjACNJukS5jViDa40bZPKDVQ5yqm7Nyw6CDPugIe7Bzb7WggXQek0VLK9DaWILXW4
TZnDaq3vi367szmi3kZ7YjA60PSNMzGte15R5L68W+hoqAVuvn6SVqFszn4M7e2BCzVtDWehCCMf
nMveMLXJ/BRLk/+8mKEK70A7oPrnW7b0+8buZRH1JVXGn6zkZmpOQMN+8J/f+BnGgviYFzFYxykO
tbDDJ0RBvjiF72OrwIXJN/WZ4+LNZCyynpwI6BQuyu2/3v3I6RbEnVPZBLoiy4prKwiq3UoKj7Un
vVGlEN2agJooMpckaP5ulPhIiTYeLs9nFcZQ2mnsbxPUuuNLin7TPrMBWB3V6aB9zeCpJKSgYsRr
MrMOC9neMgVREzUgui9kL0IyKxxPuFoO/2aL8F9YN6C5HUX8+Ur/GUrQZo04Iy5152uaMojEgdiv
P6pcHeMsJ7/j2L5r8Rp/hdqlO3sO++5/xoMdMU1G0D5Dlaie729zjJo3qPGbhyvBe644YMeJKztn
kf+MIBJc5SAMd9i9Nkw6eXqDnLYwk2dbZecte+xzs5fcE4GBRfts3bzmxPkCbucjJf26YFI9ygFW
MErDjtFabJLzynfLrxc5jl8rytyHnhNQ91/k9fBOnIyOOXOEO3YJ6pLkvD678oddVkAsOwDGiAqb
hJiESkfVkSepCwadGVhZ4+ltfs7c2QFpnTmSO9KavQsWMYmNjzfrmydHJ7jUTsUxi1NVfpv+0lwl
Yl7QouZhSI4FWkuUzMNBumuyjij5L9W1N62LbBc6vdGeTGD+yvDnMZyWqJH/DqHy8ps1IXydYEqz
WF+DexFLusewoqjrKJcbnAPJS3I4OSr3hnsMCthfK4sVpr2cMsD5YumyxfWn8GE72YNHpmUPLIbR
qnnFR6Qo8YSLtLUciAWJGkPq4ofpSvLryJg5yMycM+Arsg1pbVaRgg+teE9hVFffmyRrBZBpqoaf
MUvqigMMpKCVOanjDBN7Qb+NVCwG28Hlb1foDMBD2toXpqE/85X5SirEiCpofov5HYc6FbYVTd9r
i2Y4lAdNk0hCElq83TYJA3IiL5k+LuPzKMpdbw1TMrLUJYmE65+D/8d12N5HHUrseg1AqH838dk/
dudcyZ1WEsThtv4Mo+WBhRqtpcM0kJcliNpxJch8qBu19UwtZ7HKGRrzeOeZycM1nfjnF+aoFFTb
xKrz+cvv/SbaCgfoi4cFafZ5sR09rlvAiyShp4DxGjXrgZvzk25arn/mz/tq1tNPIaEvotyHjZQG
NgaqM83uIZlaAHzYvxjRHmr5CGdUxH5c29pzkotVUG4e12J9AYvvi3hkv705x9jknSwbYumo0B1v
DIp2IvRfoT5BrMzIBAjJygJtS3DIGFKrXowXwrcbDXqchjVoA4tpjZ2mqgJMUjeGBrCwQGgGm/1K
ZhHaemtq1IlIdUq2XyX72yft8NOEq1GqW1myHZiRKZyTzimdrlSXIuIw07u2Y4u1vOldOXcPZFIK
lItspPybNGG8bzzAI0w/vFBi583iAKQcKHgDq1CiFyHpccs5e5HpTfi1DVO3hYM8S5TzmamyWwhr
6YVTXyHX5+ckiAuEJoosVUf1SYZyfjcsmkB0nxcQAky+kxUtQcIBnGf/P7PzLLCGHoqAXH8TI9n7
5uxKzgVTK3wfNAFKoyfjGkQSo8tE2e8gLL9bTTdJApbMxd7QUuTLwYPLmW6Eu3ljg3ytIkLqJj/r
s7yPZ+9SsKHyb4STS62aVA2R+hEAXBO38/Yu+FwS+Iz8FY8s5qbyoNXzMfkk49JwOxEhtyLdn3ll
BX0e50PnH+gmvqHkG30v5+AHwiIUtls/U7yt5rjK+lYXCoSC3CL9xBYX8WB/rQcDFwXuz8SHyJ3r
JvM0FB+lRO1PDhbuLMNhpJwuILX7rZrAee3Z81cZ2MJkGo/MPrIukdOLgCfGG+uH4E0ks0vLK3va
0ajidpVt0lMesCI1cSM/B/EFEE+0kBsdkNBlWVk53StV9z6WQSjdlKzz//a6VspcLf91uLiZGjSr
xqK+/KHWnsCrUJEmy62HOM731KHmp/AuwZM1jQ73VLrnLWegOLgd0j8IwD3RuBXukSC/4mLphOBm
zYHiXztPodrJSetNjkjytr1a4QyqbRt+EmJuqDEZFdxpwcDXGD3hvwufwmUPfr350mjQN2IGA0Ys
yXa0Ye6c4wsvvPXwafGKO7WFZcNbYeyB8d+dE43cBldvZEo0maGr5Hp5Ye9FtknuRgomReaLAVAs
7LcIe6VFSuFcFoMSh1BU4I50CekcWCCXH4/vEREF+N26PZzRy/XYDkBaMqjFnvYJoYjJcUN+CVmu
nJqpaho3KdEccVoESpdg0aio7lw8qoXThkcioiO/6jV/D3wzp2dtORz89PxQxxT5JxeNurhOnoq6
q7RZQqZzoCxxCB1DWN3J4D8Hou9S4JsVT05iKvrraza8Nv239zcKL8iMobUOTQh94M5bT8EUB60g
8y5w6y/GKfDZ2K+kzYNHGDAlpNBJNoxAZmQRFEQkVXkBRkSGWm8pfC3jAl5d4+ckLFY2nLLPN31s
M2mgtKP+G08+cn1uD38NtuGqGVv1b3xgwx01zs+BxxQo7FRPVQzzhZb0KCluOX5ZChSB47S/yvQ8
gFi9R8gvvKPu5PNQghTJS2ZqrzcgO3NHR8qD3/YfZIwF6uEuGFENjNgHBvCTlZv6pXyLAjLfDI2T
uMXtYXWeCgPdH8avyZLpLgCr3XGXjSvwnqYen7CgZKvdFfVmBoVMRK58nsRNMKUv3pYucVWubcpJ
49IiTpMn9jo80Ia7TT/YL5P96lBh8fNmvMS+GbdmnDOVsdDNygsJ16eGEGQisKN3U8wX4hQhK4PI
hGpLfoVOOxKS3MCe4TF3B8DN6jJYpHwVCdzlXE9VebpiNi8T1nA2Jc37bEUk9ZjrjRqcuyfL/7A2
TpH/Wb4NavO1j3xkxKwbKoMLxt9oQ0wMkXxAETEACGagbzBL9agy4tW4m9RkckVzAmEhUQIkEjri
lLWcvk+SMwa1ew35UYzyWNoMaf0KA6FQbLB5D9MDnzrHSTD1LOqTeRGLiGcOQrJpkcngCg6T2+kD
AhFFi2xJ/xaa1u0h2upJWvrPNIcDvMUYynvLMnQSfXPOdcNc3AwsWQWpJ7UOGOrsCYAK/FTB+xee
L9aNGof61o7Z78IsN0aXw1BRPoiIEdMkOt7fvqwdLfybzGMGgDamYfDFGbI5DXfhYVpxj5np84lP
O0C7MqKHZNjlYcBgDpT7jtXzGNFMudUQik7nB4nwIjdguL8VAl4oGzs/Afnm+1PV3fDV2CczXcwV
NvnIrgSDEIBxcFRqKPmJOr6cPd8JyDB5V2Irh8+HwoRDVf5pLM7g0rGHnROiWtstbXQGWOTLAP6g
k1c0+Dg+9uPVHLubKKQjZf10OU0ttC36i09rO7BUu+3LI2OgDuV3Ma5DLca6V7PJ/XQ6OpS7YO1R
jtNfi4ZUds9EJxD0dsAh6uHjZBecvN0NNzoJez19aZ81+PddKiBNmnVzSfdVLZ0KI5xggXFbXgH/
ElXPwO/GNKwZbMMkzVHL507NdL5cADfb+giykH1G+jzHyaK56aerkW9QmnrH11EE/bbqgJq6d5vV
qSQVwQfTAtYmk3u5KilQ3Oa1sZk0fWzayug+WmWTaH9nkE5Y9RUB1shPqJ+k6+dHQK5Ak1UISj3G
ACOL/2iyxYL8LOA84woEwFlD9vhkxtUFTqGnEQtnYAowfnib79B8skDUeGsDHhQ8pwG8870UL7so
PsOb4hpbWN0q6of/W8R13QBxLu9k8L1P9lvw4F3/yva+GFDG4B67QeDPY3T4yf9cEhmbJ5B6C+Mb
457NRLg9WN/ILVwMTeVGd/Vxcs7UzVVKDVFQ9tzm8JLayRjZNouXnuxISBt262ONZyhFJh5YYFXB
0qxKtRBqwHOlC6eUFq43W6jPHfDKBw8sHTmaMBIqVtutxjuXQ4tCSo2TYOMvvvG1ClG/aqZimfH5
CRGkyQSghGtBnG9PpTzhK8E17IgSzu1FsbhVeFe5rCLjTWh3o4Xy2PzL3hx1tX8rgHU3IcuQhsSR
QSdrhTQEbW2ArePRI+MhHo2S5NwTtXzUKqCbvBzaBIoZ0RBEqDuRTs7uLKNsOHdQyd63TVCIKD+q
nk1tdXmkqxQ+GkJKvk99MFdYjgNjSogAMgXZepNtE2tajep7N7miUwqu1zk9T8+1sG0K+MYEhJl/
TxaC8gcJgmx4Abp9xMKL+HCWRx2xL/Qiebd1T3QiG7b6fmJK3bNG9s8OowSga3zFDY0Cpi0iNm4i
+x9DeqeG8IdorpasdWV2OKf/FKAzRdZffXrapK+jNv/CcY5zO+x/j1arHFoP0b5DQ++nxcN5eZOR
/vE3Vsdd5rEtoS3P+DN5sPaMMRYU5PtgJ2H35jGfHJ1ZrFuaKTxmxniKE5B1QfqLG0K4dk6mdwLR
5gyuXoWlelax6V4nA6WPRvpzQCkyLcpDvt/uUhqrSmZ64HAfdWbFaFW3ScKb0eRuK2pFYm3Hcftk
dDa826xGMUdVGJx36gc8leZ4BRPBz5H0rTix/3QmGCAZ2Gr/2m6zXS607OiJfvgYlATUveG0vOMh
w/iXb7xkEhvMqDcHI2hr73guuLrCKs8W2LAqFALrYa+SmL4/x5mRH18fpXx5bl1HHRIoEbM75Usl
EXwCvjAQYgThBGF1hs8uvZG7OWSEp+iNTtBdSwZSKQXtfrGRfUHWqPDqXu5m56npivsZIwtf7tjS
r4+9i4WqApHrwlp9BUYclnr/bjBhJCrgkHhFIT1a+XigSSRNnvpSlqNKpkbI9xzzucv6ZGRuMnUP
phX2LQenf+hfdKD/LCgtG2jGB58E4tATDUAR5njhqgTEfReAjtvJId7WQTFrLwWfE1jezcZmchGE
ui1cwnrQ/mrob8SMpVf4r9HjimFJxNenQwHYiFhkXYdmpGmgmv1lxs7wCkx7J36cFV0lA34N45bl
aVs7s7fyLr/yyJnyYBqGTNtqzs2z0Autugiw1zlzM7P8YHYUu1QRkuCyg7B0ldzZWwhmM4PtjaKg
veX6KHXWAblWifidwvhOq77DSROd+LVYDchUVfrM1/prRYirRkErDYgq6NgNfMiObCAnQbDlWkV+
MVcv17CI44Rx8nIKK6HEKLmI0QYoXISpeOdi/AShRXs9IsA1IwfeZ8vqVBSprOUzhO+uRzyEc3o8
WJomVBB/lviiWU3APLdwFqpEFHLRbUl3Xi2nsBDe+I1n3Ot5Uo+6ae53QgHaaFJ19gL1KB/qZb/E
pf4vpHt6Aw5LKtsYRtI4G9HORaKU96jxcw55n+jShERfvdQed76NdLCDuCwfGEo5lNE8fxNWJs5x
KZ8jqJs57AbwSkKSO4327TyrRiQtSEIoAri/bPYEufNSBgxKaYRHL1bBLwo5d0js8dJyVg0Ez0hv
kIl39pNK1gBV/4veACJuSWjiqPnTmfBXUIk3eDFx86/eIVeQgIcQ0jsyff7UKh9U8Yo93qshK9du
zNG4ZkVMARIvjAZVgk0OPTlCu2jK6riwVRiMG1wxymIGjSpC4dGTPrwGSh5aUi6e4xKIQQ/UaJoE
6OpA/tpfApkKs6G5+YTrI0sfDh088S5OH9rISDw+pAU+Fk6P03m/1SpvnuBF7vHQSb0JAlP6WVWf
fjnUhQamB/4k6NVZSlPDEfc6hEx+8zFBl/BXhpwt4j86OIym5EaEz2v6Km1t9GVTN88005EO7udY
TAb0PaXKu8eukKQsNv2qrdvnOlFnX8y778qdTo7nxAAMSfKtkvUul4DK1VM2mgCtD79JKzQV4h4Y
MD/1F7HJDqbgWO6jrY0FArUdnHhQ/RRPYFVCdmoMO+ynqgDFGSlyhvNgG28EeQ9yoVC1yFUyXd7/
taOkDmnWhDaBevxpzz2DnkOYdDg4IitvGYkC62tCfuPUoIpgtznPMi2tsNWzJbpCMxtX+OmbinZM
NWTNLvT3UK4I9LGP6vc/0X+lULeG/Fxl+7zxVlp/N2YbBLUmhwUziBf4hJ0L+CXSu+02ALX0b30H
6EwV2Xw3dI2B/LBzayKP3ltVJKKyU3ywjiOQ2MfmwWYYcZySfuRyJo3pL5IEOlsAGDCutQtpDbXK
zopH0WO3iebzKvJ88bj8V5wSRVayG97sqkInecStx0lKIqsw2TYMMgKRnR+MgCYZVsJarVrmgo1R
G3EqKrkp941GWkUY+IZcMAyvQJJDZEj9Ftyio2WfUHV/B7W5yqiDWQuYCe5B8SJNZT2KDv7DhmPb
moxiR+IRNoQjF7ezzVQ0nDp6h1hveBvnYzwxTvKAPJ4vKC37bdpDOEe+k1CyVybXXi5M01OZUAJZ
gC4KqJXC/iVOinzcABvyHhS+qkezMs35CJxQ67U5WJWsSa2HLwA9uOIXMwHvtyNbBiAaLoYKeeE2
bRJkUGCDnnybqjdzcNB/oWhJIiJ+Tw4vUY4Yc2T5UK3ux0DSf7iYEYhaktrZsqA8RlA4hK5qdyzs
rQpbvaQVB8WcCKIfoO4mnzUP58B7ZHYg/iiV0HHKA66FFney0Rc6MfpD/XaBTHRyz7KSxqBnwfi5
fPB9MmIuZymlCLa05IW+0+8FQVIK1wfp6fD7L0VFHx/w83t9lS/mgIXvFMwxymSTVJihYOJNmWXf
qNAOkfaH4e+WVhzQKIccwnVznLC0sVjSBVKGxDpUQloJK2vwpGjxvkjQcmtW0m4+GgxK8gDaDBnp
E1Ys4w7UBDkBTWI1csEZUbdW4mib+i1o39+/mO5ZoNWBQAUVwShDQZ5fucdUJ+YU3xsD66PvWodM
PBGv3tCdb7qbSXdadIadzrvIekPz6Jfb2Gv+eF8tWSU47nAWpA0j0vQ/V3ONWqtXKcE693fjX2uW
xTH5hhrz2zGRQ6lI2YP3011v/SMKX1KtGXeXZo1fXeUKYC2ijioxtRpluIQZso3BvWcOCkFI2Nip
1pvXb/yEhjzJDU7vFqzKLX4M/gJOSWiAbbw+HbJcfsieDAIxaybPAg1PCLzWyXM6BPftojk2DytC
7+RFuq0n43EWS/JWxFG6qsiYNkW2HltjLSk4ekGdtsVxzBu9DVgi/hpWL6ts5cVUAj+cEZPc3g==
`pragma protect end_protected
