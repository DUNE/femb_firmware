// (C) 2001-2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
D5JRwTjzoKsPqY3eNg5FZsmAz1uyiU79+bp+TNeOCUuvjqATiRTFEditO9Y/JY1flvQOuO1vyCdA
cUIzTpU7uSp9KH9eDAufdqGF/CCuRRCluNW/GLjd0GpSR6+pgNBAwnXKeenJFLh7/3LUFWZf4MSC
uXkm/HRMHMCyF1qwyPUI0AEVInuEDC1O5+Ocu4lw+NX+7yrMa0XK/1L5+EJ1C7yxNiG2uHtIt9zD
2jllki40e1amK7XlHEfuAqAvquhlpgFh3RAyyq0OHxus2u51LdwDu4FhQrbUZvUzj0Jf/xNrLpgz
zlfMenvc3owsTSYQtX2KbyuYOIDktxukisRkZw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9456)
Jv/zHMOVyHhRc3sVxWPsOhcUExQW2FZ5LFMVDsWyPR7Krqe0BFRZJFLma1IlUTufazJ5+HdmBGAS
5daGMpepvSVbyeva11oo6JDPqSc/j6qXJ7dmd6GeU0z1eWoJxHj9eC9hbilPeowq//fT2Rbrb/d1
FTorXpCKFcBvk8ZQpr2DssB3w3YGVQSMiQ1BH2Jabv8vkFBKetZjDY9yu9STU3VRd26BITuufZzi
DVZN2F+E6h/5MV07hxVl7U7V3JXzk0zFxqrLcQ90rJgDMfK2DvQPxHAIDS/rmYgt075LIM6Xtyjz
4VmSi87Qsz1qewRnRBTgaW9szLsUQLxQ/cx/dg7Axa4W6ElHM/VCUYOuRpJ3jHWL+yu3O2oSZ84q
ZqZJ01vmT8u0tI0Mi4EGLgvUbqvhJyPt9Pb50wgQCZkvi+TmmSJ6dmGBYH/cI3y0SRUTkJtHWew7
H4VKR6H4Nhf4eH3yINZAVO+VKg6G7FuxJT5VuovPXn1Zm9a3HhnJCW3xp/9KSM4U3JNMd24u5YAv
aqJ58RiGx/OGSWKF/M0aQp7zNrpfrFc8CJGWGlOb+WdmM7k/aVbUTl0lZ/9SFYs5wVphz2dg4X4f
QUuhtY60gRa6iltKRoBpB7b0fn6GOvMkkCicjYVqTGoBCUxtrJCjRQurFfyhZZl7PyIC1+9mFNep
6p89xToKCfHR7f8U9ckKaPqi/9uhU3zsCEouUFO0GS27uO2JxEGU48/D94vIDeXrK/IezDKqkKwD
DvkowdM5rNhox2nmOsIEiqHHolSMytmHnO0fNXCozGL3YLdMqQLiyh5xgi5xACUGUu/jKZvGvRC9
VtE8p+VwX6xPN5mwJLdjAranb+SdRS8XeqT3nvqZyAsViOr4hnomnESk8XY6QGHLeYFGnVixKPyG
bcQH8CE/ddBkutuakREIgTPMGgWjJlapaO3jeJtQWI59aS5jYl2ADxTPqztJlyh/nBgmYdy26BK0
gTt5roRLXMaY/T4cBAisEjf1vhQYkLat2NK6MGdVFZ8uUiseW7hFwyJJAhfJLoMDoXha93zXIz+z
uz0IBywq3nwFJ9bW/sAQmEyCDI8vQtSNkmniCd9QnyLXUq0Zcm0nKi/GotfRN9pXyLP/PEtrgA+E
J70s1DBFfF39DrolgpgSnYOoO3vyQT5YOTBTeBcghodtWKk1gb2rM/dz1ylPqZfaKDanNdVgnlqd
+Hq4jtFI+Edc2zKvHSlmLBTalNsDDM6GdqqAD/ZQ1Ps/xYou87dDWaGqUvDF7zvP7sx1rPaaGyRN
9KFQ4BzZWBXBD6m4FsbygUe1fgtdq2/+EaYUvp/PoF1CeUO1rqd1svlJPoJst/SGtugDZxlqyFME
QYRig4ASwb+Vj01YDBhS2aPPkhM4G12T4Zw+c81cIJZmEvhHqmIVOeDgRCrf3yzWga5FgxNDZQwz
/EuqDTRiYt0Jh/ISmOqWiS3KDrZbqiY+CJ8UZyQ/1aRTJ/YV0GVvXaaseGeq7QdvzXBLVwUkB/FK
M6pHsAnxNPTd2jaGJ/N7rSbS/9EqDTtxImwUe80Lgai3Ubmjk0BbDBvCJd8w+k3wbyCh2UX5eAfl
GiGU1y5LApCBzMWFVGwn0Knc+B+VbOdk8b4ZDiIqL7z4oSkMq1vMwT2NkTibYkYj4LyV8YOCQR2f
i+uINlzj1XkdWM5S24ZiL/a+GR1775uNxx8q6fMBvOU/5pHqZToRIcDJspYRWnULIF/6yHHZxVWN
7qxljewe25DyetNJ6dbFS0TiV6manQ/zgZHutVmYZ/nBmflWqpT1k9Us1acaIwArBGOLfcoCd6ZX
FofwwU+SUXI0eraCzfsWxfngFeSne4EAIrCDXg2igmgEzC2h8qSzzNOriHSDz4KqJfLPQvFBXKBN
ClJM9tdYAqOp9YktJyYPFUrXXnmedhZPF1/uzYuRlCkDbIvqWhcr3C2EBb6Zi7iLRQ+rzrdNFs6k
pMZSaNk4EIwmj8jYQkkb7u5lZQ/K1N5iT2B3aTD2lwE2D6PT113F8ieo7PDcZmAfv2jORvXfmLGt
L+qQQfia2OckldEOZ6D5YZi8eepdXs7H+D6AtaOLk8J6jqNEEFOXT2xG9z6hZzPiIsx3KEbsDHj+
vjucH0Zo5/0nMx3PSrN3N9lZpzqjTVJcBVl9ozEMx1VZzz9JLnbWBgDSbJTbmNnIFGFFRUtC6f2T
Usa9ukL3FGiCNpDgOMq/VlDWDHHwji9v+0wxZryT6oVzQhGLf2jtwtUS7f8QelXQyxs2gzrbw5vl
HsXTJ4M5rFNIzIRQvvhO6llUb59k72PWoiEICTJvMPzamKiE27nyKbRr9+XFuCXkvay66SQTRH2z
28/6cGBTjvrx6qgPDxwtgv77ntB9C+aU4ZgbqhOMob5FBKCHgnQNuwIX5kqW8AXemmnjBWbetQAf
lzMXhkOFPsu4OnCxfGB4leagmAk1vkt72MTiBWvh+p2HaOKTGbYV0NziAgB53kD3tURgW81GT8UM
Gx0/U6pQidHuGK2T/YlI7k4X+4Mkw0pKyPlBtR5XdEEFXGSxcEILv7cYIuxRIIMrBhnkAH6HRTuq
FmKq4iednLshde3lDw3zI09Lkv2D8Zmj7Y586eIOyWvH3FKs6HdYKyeQs0B6DYR9HVu0ht2PQRU+
YMFOrlUKsZssArYFY5mnAQgErflKmEZBwGDseP2DfVG+ulXgPcraar67oMLbcB6rzTmkQEgzYrbN
KOdwkeloij3r3dk7VBWxq6jFYKfW+5iUx9QqVjU+AXH45hHHRE/xROFodjgmmwrRebCLSANwNnc4
IokTggR+oX19/KoOJmFmVRcrthGD9dVUHAc/LWRojLza7jiNO/E434HNCe6lNhIBJ9kzwGJVzQ8q
olib97YaaNedgZHCfQV7QKQ9QKxr6R4oLbiX7I1AqcVhK9sTjm0rTKQ45xXLr8xvxmUBqjBP19mb
g/jWub312FhJjFO9+ub0oml+CwBPLWWSM9t+YnQAv7SS6tYYHwWkCeNKQWxdeAmLUV820aeeMEVP
M9ZuBVD1+T/S9QHk0IgR6ksNePm8jrvkaFa9QwprRLWQ15tDIWvls9EXwz+h1eabaLbDeU2++0wx
3AckOeCKMVdoZBeEsnahWDl+aS3KPSSCgwfvb6ZDpE5oJu1NO8jg2p5RsZB6R+JfA5dXcH8yPyjT
28WUNEbdtr50yaUhW92N16NY9aUvb4DT6It95kRWigUiPeoNLZzZ/E9UyqCrai4FvtsY+OtG78Gv
gtZM1YVaGiyx1akgzcRmdkSrJ0OiiOzWGOw08T4KrrirVYfifi8TXR4gTQxcIykNHCWd8zcCgZ7O
okgEp+VidQl1JB+IfJsYEvdjquo/J4uJT5LEIaJfQdRk9QYT2uzCP92FDTwO4McernlnIitvMP0N
wnG5vf8//ufrUHqb0sN2QPIqAc7KWld85Af22c6pDbwlhf2h2IWQbl1qC2y6itjqq7AWtXyBbue4
sjtH/ZZrnljGFmfa87GQKXmU51mu2kbFmArIQkNEbG49oY/Xd7Alhy7B24mAQrEFBx/b4NWeX++B
Z9mRDC34G+uYulwVbrxij+PkSnVaVwY74ULb65XemED2cCyYtayD060h54f5BS3nrF4GyL4USYBc
LWBygX4zBbGRpenMulZ71ZaI+p+BEchC6gjOQOKCcWeDWSrcPz/B0gpYuXfLBfZ5YrtBO1XbeII6
nS8rhFpC0A6lQ19kpwb9A0JpYSWkm2sY7Ee1MEec1jgELf2jlTAxr+AOzG3wKbHwBWHJUwOwKxTY
p9T3zqIuPpOrKLy2wb56BDsMxJ+bajhkBoMQaD00lTrt1EfNHntzq7JiLBRWM+ET4vizguhRxTUe
bui34Ik2PBp9Bn55kysqEmYlJX3cmQcwaMe3P+5jJEYqMB59axrEFzL4XleDMUxZcfxL++prdq/g
dfU2ocIqAAE4Jz5BghoVp4pudM32ZyOuYlokThdcMkMvykCFa5EId5djU9wjY3TUptDWvXbDb/Dg
7n210oozP9OGrdAYp0AOwHnk6jlranHKjFPvavug6fCKSI8P6sLal4dwbPCiNTbA0AETl1Md6+z5
IfP8SbRzivr2VxlUM5AFWz+ZEP2/Q/+XUPvXk6hyvZLhheLDmk3H1nTGOYMtRudowXo5AYeuMFDq
LGA5tlLbdToVyLdjpr28DfD/E5DJemJL7fPGLeswL+/wvK99gTlacjgccDwlbiyQ9myedNttRYOc
64azt5vSi5BMBaUHqr2pMv26IivTuAvetbqxFoIDK+fU/SmLK4/2oh+A+FOMW8LR+tuG75WdtaHn
W4+q1dbMbzEF6GjDp2VRNi6O3EbcyyG9GP7BfCtBveYlupkxyRfMZ/wpYgRYEyjAx4/soY3yRXLj
+pi5BmjcFUwQAAUgOd/30OWzE2hvKCN4PuXhOTEGK+sY/hpCPsHipzWVcx6bDcScG6FTCOUQ4Op5
4l/Db27BpGYCgikQmo0+c3s1PpyqvnGIpWJ9GzDxhom9UjuJiXvyrCkMQpqOdHVGlCpUz3mSBmnT
cGIXYF0/ai57fSqE3J8rWLgsH3YQMSspk6uBt8QwiW+xYqBnV1tGkt/aVL2d68OIOtIFFdE+lpY3
q+8y8Bg93wLutwLprf1A/9RTrlt7/jd3CYlmIOiHNG4uGUd8sUWx9lYGTaChvlqNUJmOp4hWxW+I
HKyGZKB+BoHmfKIiRgaSY4vmix+2S8ChGJOg/PyAqlov/6hIBhIqFK5j5PesqDwWZaEpf1H1OliU
VQ5xRQQn4jRxvSWyf+HIg2yPngxkRv0qUiKXBFweaIlj8/QaTrXwkIBwyzSzRd4xzkE39k7ZXMWd
doZ7lFomN6n78/yEcHsmmCxBQ2+TRxdREEtO5YwI8pwRTC+tiI1V5mRfDDTze0uqDDTDOlImAyV+
8TGCNCfR3EtV9hyp8KfPHeSvImScI+45fNjHw/SR8qDzLU2B8HifZ9bKctz+bPTGHse55WM2QeZK
g6q8yPvP2mr2JuJV/O41wxODpi2UcnzR2DohMG10uro4mB6iPiWrVKVfhPMD/gWebytfzisFi0ap
9y7jYE1B763LuVuO4kU+7hBeQUcvXIOTIfiCtK8CneAVEOSLHZYwcexV0Ktvb/mp0wiWJSitwdhG
C6EcsFpkzgUB9G50bIj5Qz1lh5qzI49gXTM/j8Bf4CFgfaapVS2GjJsbfTfQmYf3zcgkAPKelHtH
S3mwFaW1hkS9KjPbAoJ5dTkjkUkDonL5IFShLyXkyPhBMP9C5ALA/8MO2wmfvHFIlhTSkyFSA4PH
xPhf5zXc3XjhhFpg6i9Djf8y5u3sPh6vRIBv41m8/tqHMqoxTsS5MPy33Qk2EEhn7A9te19ecmPN
RPSzNDqptfzjOwwQGc2m3/0j9TA+WYEHu5pWeSckm4WyLTN/hfocgts9yZKHkZ4+NZgsZ7Mnx4/h
ti6N1IEgjspvXajKt78VuqZmDS49K/+46osYaUDw6cD+a8SGoJTgl7hs60d0gFTatRza9ftHeJHE
SoJvBPaQDuVNdW/6KlGDttEdCu3C8TsvLXgoveuLSy/ZZmo5dO8ca2vP3zy1wq3JxbaHHtqWcQt4
/8iKxCLXMzaIWI/y5wxAu2llOWt81A4Xxf70NW9BBGuRYkbeL/oHI4kiVBKqc/b4qumHy50KY1Hx
GYpZbjTIoHIYnkiywDrq8BenV1DRyju72Cmw1PTPkbjd9J7rdeFOT2BP+amXW5lYkpCdqTwl+rob
q68beA3PoymW4ltP5bfYOassQ/Bwwas2aup4rsEcuaAbVMZW3y4NcZq+R9EYK9oAbQ76npOQ5cY3
slR27Crh7GnQZsnKOlqKe7y93h4aUNAWUBq1toS5ZzcROEFMLSG05n2pZddFE3bkpqDx9FyWt2sv
cgvYb0nMpXPN9q1g3W9gAkA2hQSyTjzuluBSh3GV7KM88LZqYZbbcJyYdtU/+CZsXPTgfdAYAEET
GBjpMNCR7mq5Z2e2PbcBHHBwusuJG1mi/NDdzXBmZEVYQ8i5dL0cr2XJ2mp9KGVfR+v+yAm4kk2w
WkwdwS8TfmgHqalK8aoIdvbnE8Hgz8kSIkpxRQACcc3+DtNzJ4t7lO+S1zHuwMpo2UiCBohylQ8d
Viq2GLvKDWCzIFUyDOlXMa+H7YtjjQUd4YeyTud7juxQzcB2NU5dod0J99Io7Xg4cHbeeJyYHDpp
FC+d+hRy8GT6sWX8y5NWcYWDCVetHErb4qCreZ687BuEBl9yzxy9qEswOyQQGx9rkWpBqTx4QUc6
7YhSDcfI6Y2Y0hQkpOCXfqR+dUBsYXvphl17piwac2RruQ5xLaVMiS3ArsRCYfDs8cliSSWDJX3+
yC70YDw0VPSWjbRK+j9Ay5zZGJ99imzavfpUNcG3ihk32dm597H6OXxMtn8Phg73klmwaxhroJTs
OPTwDILZoGo4S3oCjK+k+pAFIKtbMrzyR9Ny2AN9qZo3x4BftNU18dMVs2rTyWYhbPu+5EJARMNR
ouTKFuYqiCfXpX2pi4UnuNhVVI775dy/EPOxvaHcfyurUGd+JnL7OEt1HVFSNeYLeADLEgQEJgOK
kk7lAVMQAKrAStJEpGJhIiTzyy1CmFPeW7HazjberN+84iZC5fJ1efS4LCpdGszAbTVnUBmc1GI3
AZ175bWwRdtnOXKrF4YTpfWWsBxYsnPsu7YzO+mn1GCrcP6EvWXLTBXUTByKhbVFk/gA1mJH8lc3
6LQTNsNiyPAtR5j+SA0OZy7Ti9ZzVolOr/r/aFGwC2mwo695GyDAXEzoRClQor7yZnQUAxFzSoXE
UY8GVjk1VvQxf7kKieS58LbrxaqpI1NXmdIRDnV2ZEsTGa7H6rTEG2a90fVXJxXMwb6LFIUBwbDJ
G0EbKHZUURyGQJ9RxPA98f1Cy3BhAc8EmnHSb/c8M7D1XBVkP8FbXRh2zDn3/aLHk2GKI+EaysEH
veCpjDzSCo7Ub31e4pBsnkBFFPW2vSM6vvUg+MTC1QYcD9wqytvbD2XvNuR81U6rGgumZV3YYi5T
KybUQzqQM5NkDTWC9PzlK1Q4wK5pM2fK/9xNKjWm12JJR9BTnEU3sZrsDPNIJxOLHdKugFQLstiK
1nVhi3xn/639e0nYge+AMNMLUE6bYxvl7NF3BDR2c99t9nuoEYfozL84eNM1tzPzgzllJu8sJs5d
w82JzIrKxV9ZnUgHnc1nWf+qlOnNmIrhGj0u3HL8SxB7vvLwJnT2qcVkhpE6VoOXwFA+zwH2A96T
eHZLF1x1H14vQm5Y0jSxc4m6PtlSm4sdTaDOtWCKQGVTY48xfHB3IgesXFWcuJAGbc9Joylze+Mt
sjIk1wd506YGlB/kfKPMnWFhDJVMQJfd1iRTR7Sdx1SYsUKgG67kJIMda8mutNNZoSUV/L3alUqg
YpjptZnTevmcq9pAJr+D7G0r3QH0Smqb00lfAg8kLc6+V5g1hPbic1MIJ4+sj89keb+LmdFZpTtG
u7XXgsIZXEljNeSm4F10Lp1Gz+dIgdLxRlFgYbfHI07L8FRCbbYyfb2QQJevnz5kQaNLWj+P2/vy
7D4W09TurefhxYDpoI+Fmy04HaUvAl73eRe0LoQW3s0tBoxtfl5TxO1f9o2yyBKCQUvDqvm/IeLp
2v4tQ/hMzVt8bBM7scw1+6KnbOZmmP39zRvAfXy7zlgfZlIg1IGKMuXVa7GRPeUOuDyylCU3QxX/
5TgODu8D2hZZTlIImoe358vyF1mg90bYbvJN4wNFtwnsaQRZPC7WeyjhmTJkTz2aggNEJKY7GfB1
LiBHSjFWtxUPJvVCyp/V/5F59MKGGWWAmzdRVqvh3263njOEumK5Wu+fcOqC9jgAGCEJ8OwFjuVB
jQL5t4dpQZUQQbZiPH21ES3N5Xr63y4LY/DiaR0VRYG7UWzzF9d4F+egZ7nRv5HV7k+Jd2Pvuavu
iukAYXKOCpWloHk1wOmTUzqKxXOhahTVe+lY8HI1z+NohswD8Voh/8lT2VgVhEiiUb1hkZlugCPr
FULdTL/V0ZiIxjg4KNfjVII8SXs1FBc/TZN/2+TiXk33OMNkExXTYPO/cTEXs3RAPhgxddOttOYI
WSsHKMRaAHDtRL8HPhgBjFJh5vWgrnSi474RPTIGPCcPZQkvRkLbrEDvrVhC1uNllZgjWmGttisW
shfcE49l90gqHYFPkNb8Clzq5kndmUVSmsY6GK0p6n4slqwxDtJnUzUG/Ap84QzvZ5I8Plxr9oas
EueJN+UfcPtIKQCbYLbvi1eo7MTGNc2SLf7eo0lFhfna9yTrCsZ6s4F79+TrbhfC62Dt6WNQtWUh
+Y8ynlxnj80yzxF7Th0ulwHeIYeHQQrbC8RIPfIpCRDr6gSqNadlwX3L2QQB7cOebLVD8Jh5XEXJ
r5+thLfABZwUGTPo8uTnjtPUz2e9b+UfyN+BYraK9N4UoIi8SdWKnXaASUXCpP0Ui/eIXD6ru2a1
yBwzi/MfRLu1x9TyTJ//eJl7zX0Lv3pxOHZS86C6rG/6PyDgZF3dzYCHKd1lgJ+2cq5e5Ee5M6DG
3c4kPFL/+Tc6DjQwqFP3X2B+zYArVyxvfUb/vSblZ6x1Y0/f7SfgAq3aK7KXF4yZXxwSXKFs9oPJ
zEkDyQxXYZQ3vJ0AS0CCBbA/tpLJN4QqRsSY+znLasq0RYZZbxqZy/LuvRQprdvIOR3f8PhYTqdA
OSEcNnoq3uUEGstiAdSGQEfrMod13Kpm2hr3bva2O0+jswhHirj6ZiNpWz3FwXA+ZTCb2hhBwcQ8
0yhnNp76XO4TLIyGQnjf7VjcejU53XqkpgBIFPlK7ifQjD8a7ZZljgXCzB+hJ4QZBsOXcZa499Ds
RnbBW+d+XSxDWsaZo4umj2aUPWCKP1ig5YkbUaX/sYULucSz8v2tBbxJEekP0fFnYSx+jIfQBEyN
iTWXs9Ao3Z9jtzeZtxXgJ+nKB2cLqZk23FqYRv9M1jUK0rrQiSmmZCe4JzqBjsnGbp7kbGWjYObf
gGd7LZUNCLlojRxvnmTQixrlqUIlAkwHkUSQvPsdsgiDhcpwB0+X4YJHj4yaJeaZkEcebWxGtAwL
5XwqMUEKu6hCae2WRS6WvCzdXBCbJyAdgdQ27TW91sh9VgTMPjx4bwBtB0aTL87qoGUqdRV/bYJ0
p37KhucTtNql6veffhT4iBHSGOF4Ia60qchMzoBgG823YswPDzctlqjzVY/GdCzrDHlJHME/481T
GkoIHAWdh3Jc34j4xfk3W+f0C7B5NXri2fVDSpBLwHkrzVnGMxnB1+rXSNsNBgo171mlNSoiKAGV
KAB5lI/ieepT4a7puwV27K63g++mdAFSINOA3mayypKilsWtJF8Gc/2YLVOfrl9yA0wtXHDiu/xb
qXgpTzcOS5BcytYkoEJa0bxAB970+RZDQOQl3/2iVu035tbRZEP9A3p0i/cXVll8wY4t3oYpbPFn
mLr/uraxo0VEKVnyoAEMi+m9RjDToOoTsiWBY/Sv2gsmXzTh/pUGH6WR67DQrMaxDPjmTnEHzfjv
v+pzR9W6GarcX6UTlNe3wfIgydE85VdBgNkSABR/k0HMNE0Nw6/ehy/OQ5ZyTb5l4hi9GfTi8jwd
ITHKV3Tk+8GYqO79aHKQxH3gzl5jxwp/l1E8sC4CRnrIXfY9ne71EMwuLzfg7xZEA3JG8dpThm7B
+8tKyj/gEL8Fmrfc0HW/9TOSzEDi7BefDrdrxGPSAAg3i1djBs7+NPAPeGrvSyOuQRN2ZPb6lD6M
oDTNztARcR9Pf5lEQJlfhdsPE8Gi4u2uECIyiR8fyxrMBhYu/oYQmJBF2xCnpqxWp5oPR6+LVODo
SUvN1JTgedbh2FNXhb9zBmBCJ6AT5yHg1LERUKnlELM7+Mti3ilBXOJNIstHivYhw9rYlhT3uOHO
SjP3AG+yMl2pyEZhG9tgUvLH5jezh9Uqx9j6gCfwvnI0ddMgyR7qD5qIGFgbbB0ATv64ziMFXSWD
At9J0XwiKuM734z2MHMOpkTKq3YVxY6mZZVpvYhIjyIx7Kzsgz685NzvqH8BJ0yXEYP1KRes5gp1
Iz4/jJgfKPLRwLjdDgx3Xc4GVisOIaZ8fBcnvssChjOP92DS3ACRkzL6tKR10LLMQzhvE2QoJP+O
7ZlPSxYsEUiDJ2PRWzd6IlWlQRqLL5BNrCDm1L6DOntTFWQ1Fm6LT7+I5vcru7QMfWej4urUEpsy
4xp2oCw3xoDOhHZT+8Dbh9zXRdW9e0+EyFifm/1JP44QrxWWGGec9Qlgtkk4KWE2bv0keG7wR3R7
xsfUFasiunVJnbUVHFrgetYITITb/xu5orJUXfp07GLaj0sHrhwkOKIuYUi9DuIhtgMlWB1JAz9s
7Dl++uQk5qnRHSiDaQTOgoo60ThBNXzReNQBeJyKB0qYJWjgWHrf/CkCPz4t1+P+hlsNsqIoMPiR
hnfN8YKnF9NZhi/fnenJWt8LJL3ZGkeX9bMy56tBzKcxV/HUoaK1FCkl1jtE/vW+SIyJq0XEgviG
8SJXOCV7NVh3W4oG194CLLxcZXBJ20fN/xgvmnKHs7BB6NtPfg90omDLTkF8+rJqkk0dMR4eS6FT
6w+sHnIJP2f0qL7/ZTVF/Z1sEIPBsDdgcxy3+HKTD7cRnXoX4a3XWyM4RjyVMYiJx0nNp4XjAkV6
nwvKhn1TmEN09vQJ/MaHpemt84e0cXe1nE16uqlvOeAyoVEQv4DwQ4zaM5PRHhQ1UzVaNSF/RUOj
i/m64Y+bjunNwqE3kh1mo2vTI+BdEEl9+zt+gM/t724UEY17PJRUu8h/VrFz0ScpOiDeJ0KQ37TU
Ov4bC033ygYH3tYx5GFfZbyeS9Ejc136IvL7losFQZ/Qretbg3Y6LOvHC6qnPmzcrFc7+VGfi+YJ
2Is1VhafhslAM8hvt0thinWEmogCC0YqECHFpYhpv11++j4D6Cv5RVWFhcPTV60EJffvVJ71qi3m
qXUGbdhypj+jFPdI/hcZqIlhwqUgwPH7H2jNuCaqC3KYxiJSHfunQ5gB65xsBRyp6PjYIB3ydWSn
f4ER/R93TMOMx394eDni2Zl8bA9OQQ+15a3xzzGCbsDboceHPsP2E2gP+klvzBN8LP9XQBoqHm+M
rhN6QhBAayPJ+LT75nyI9AYmb3t+dS8tXu3wiGQq6jKDgPoKDnuVK6oAqse822nYpR2omIZ3St1M
gFYSVsnLED52aoRceP/rNm+Ncc635WpNEWaaif2nRgefYfgf12sALno1aUQQyIGZCwZPFResmKNz
4h6J3DY1Q11327bLRKJnKBWR93J53igykicNQr3PKuaoutjo3gZI6T4VC07TmYG6mRORrhitaF8n
qHELertN64Y/uSKpL2V5LTlVtEOBe9PeD4BGKDUukrM0kV4JYC7OhcFr12poKs3gtlvmGByGubdS
fwO4wLFTWj3XBoGrOQUDZu44KHQSmf6c1ljuFJiJItJ4G9xDsniPPyNILkGmD6u1YIAoWivuLn3n
Be9BDE2iBPksl8EUEWf1WUIYErKP02hFmCr0c21bv8N+Dx+MsFeQ+K28CeK0SX2U19naqM5cLRH4
r+3Yt7KvG5VJ12NhyUSHaMP29H7qsmhUhJJ9vtsUoxf65zLz1BYJ0x8I5o/vk7M7e2OVl20idvmx
Z8DpmeRn7Z4wMsKLhbnJ7F+TF6FtPHM600TG7jZYblW8ioDz/nWZF/EKAiZODTkD4E+JnLXNhwCF
6dxi8l1PbIAqUvwuUW6bYSv/9ubSLODZQM+herb0sR0MjKHrRYbFSDcyqJuxN2j3/lM1DoZ2BoEx
K63FakbLBe+DWePEaNzXtb8wmQqvmMcQLH/KzFIyidwrOu2DWIDVfMhw8+MUdLdlh/JxoRKHfZMG
kjXdOtwFPu0eSpatq2q3fH+bPOGEfmJ10lI+3NO1xG9DCUmpnElx/vON2lxn7WvsJPjNgp1Rac8M
jx3GT/FOe+YUrqhVWai+aLh4UxyrgGPqqKLdI7qH934Q1u8EhKmjoC4yNjJAbje9nqBzDt0c7Lht
Sa9yAqOeMHu6n8O4cfhDdDk90xDeXcLUpCsqT3KoRcRSyoFqGgzc//yHB5N162HR5FwBLniWmuVL
1bKSngzwPRudgJk6zEXPnFZKLw9Mq9BL6TinTOWMIpgL4Ax8K5B9fe2dy7/1E0zYxNluR/wYXC2A
7qjoDehczACb8upMR4tlBDHUyL4gwjnYs0WU3ZB/xKnUiggAmA+PLVJs3HYsux6ri9VEFE2Qp+1+
dbCLnJ95guVMLxYrpgxeeu0Oy8V9KAq4hMygk9gA2cVb2vxYeuepDVWMKldxL+CXPYIqJGnHZmDy
kJ7Y5JhWbvQvF1+Dls8x140+8u9Ej8ea2OIBb6rZ7+fed9sfk7G8jMKGSzbOH6rpw5h5cWeiffGq
DzxxfsyJ9ap4rlqS+gjmtG6GUsplt8VV/Xr/3Kl2Uw7snMyvddHqhriJ9XASMWOwqX+kUQ8wmO8a
c6hXkRjybGR14CLXNfse27NY6nM3BPmwUPj1fmy4THg/pik/U55orY0fH3wGJlatvIIY
`pragma protect end_protected
