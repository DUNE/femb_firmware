// (C) 2001-2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
QIkB3L0q0H2bUNqT6+nQB664iAp9CfWUR9E1vOTgjG/og9t/dxkfjwau3LGvt9/WJIKwQBZJXHpq
KksDFrLFp6oI1j9sEs+BFCfohuru861qRbQ66VYspVS3QZgjATtujmwJmS/+WlRiiIGhBMdoeoFL
WSw9BJ41FzSPgxhhGB2L9QJtJ7EeHSKcq2tF082SboPrUgAoZb6X1PHLTQXscpMefeChMAf5qUQN
bRUaNaNAu1KKygx5KbxeZb8z73zwnyHSZ0KutVVj0dddM/e+IJ8MJSXdjpD4LuGHEw/BOIlmEeNS
btoHJ33vCmyFVphqY6Xgirxilct59o5lW4A96Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10960)
yYf9mCz5o2jYdYf8F5PFtAr/XCACErr4uLmi817siciAwMTBj5jW3aL7xi524Z7B4+tXajBbPLt5
iwEH1+lq2T1KB7N4A6YVLRsyR99dC7PWa3W9y0ijfWwdIOPT2twhpaTVXqA8q/xcULu0zLGWTbNk
W6fdpsofCwJ/Ft7M689Pe+Tx8hL5es1Qm8hWAFDuNFkYdMwhewQqoUV+NbJfHHDKA37XXgRAzqpC
18jd09JK1KPm5PcdZ51AmfvjP+7C9ZRA3LZIkI1VyALLWpqGCCwQrOL5thF3iacfwWgzYCc34HZG
CHzweTNw+vBufkoMcLTdTO/9havAauRm1/y7ZX8esQ/iLgEElKtevhPHCpkkI/5CGVoqPz/NcmoK
Uhd/TIS6nfEogy1ONG8o+X28jOhSxRpohbTBV7A3sGaiCKF+svdxBtlAmOWwxaqY0yA9283O4VKW
H5cTW66RRxRZEU4A87I9zeYnxeTUOMAvjoTfIZskasuZ+hozMRtrDnY7QHq3g3S4fApbSUIaGysU
CxwDPZtN/2SIQaythVvq68xCnh8WLrbXtADOnvVLcHsHCQ17dRiDv1ZvkelFn8T9vr+RTUvOMipg
r414YeTqf8PK0WrTFMNSuhmiGYKX9MOv7cPPXfAVy4CIqNep7TxnZ755Z65+d/hcs1Q8YU3CHXVq
b6kIFMRpO4KwxKefPdDCUPZLiyyJwmaO5VdoXo5y8MGDQLG9qNdtUkyOgjlJ0v5Rg5bRdAxGReIA
ZtgFGFwAbYaRoTclhDyb2uhd9xJbcunQ8Ym8wHMxgqenjQ/2unCu20uqj+SYAb2ohfxqyW8A7S73
llmYyOTnz+KBASFfA/g+Q7hjSkacAo6rE0dVhAksGecRHrbMskb88FRGqpXzn77BPGPAFlWlpYQr
C8WqrklYeqobo7NY58Lz9uVYI/EmdDCo03mkYhamdPmN5zSIMG/pNtx0chISw8Kes+dd5/Iso3aH
aw4SHLuB6UF4vmTDX44Mx9jXdQxBFU8gsPsbwebyvrWSybB+z+uhQkk3LrxM7vjRzS+Bu0Y0aGnh
7Htpl3R3uMInehG+2an6DB79O1eUXKfAWzrY/bYIsDDYW38DjJcKZt/gJQwgBZ4ozqxDhf0B4HGN
/3zOv9dxbwfuEAT3HmFzDU9oTfOwnX5GWhFLCNpbuiB1SIPZLATIdNMTwR2POgw9xvcl0V+AazWN
WMhL3Ojt4O+o2pinjBtNP9B6FlEVI7WO9l2ynHBIvlotOcntlJllcTdpC2qhpQmJgis0vPKviSFR
NCS2/x2+tQWy+YzQu7efkKdsrraI6U0bXMUm6hyCNeT5JumgIaAVu5ssLcDO4jiTV3PccvCwKBZt
Bmq2Jp0wnEiv9RLgO3QWrWx2MXjm+6xYe9wo/ykeZOs+3PMaVVIbDA4x1mkIHS7jArZkt9g9TLDo
E8JOJdCuuxSprx7oeKRv/mlKprZL050gsbgQqdLGIPOvX+b+CUie9TD/uMFltpVsyHJnXneVKl/l
bv1GFx7oMjbbwjFRd4tzjMx7hRQS5uEa+xGwEedjkC2u6NUVix2g/j+0Uv2BCkGLr5uj3eTUaqVd
qbP6on/8Bjj8KSebFCyYtUhIYEjBxJ5FKfY204ynEBMpHFqP9mgeJApSd4E3ppsYkiclwEbhGlYa
QZos6RzcoYeiu4vtkePX3+HHvBxRGPilA70BxL5YnFW5hPZde4ph8PHOQbfZv7TQODzbfrDUyrXm
l1iDnen8r5BoNQ9pDgkqC2wC0Jvd7vmjJKNl5uJPOemoLcRUP4DaZSF+0a8dQYoyipvQod/Tn64Z
7pG8lRDVn4hoLxeAARRxom1XH4esq1qz6qRFTgSqBZ5+3cMf94wbeB/uqu0UDoMBQ0Y8MSKMTQon
vwOD3FDDzSQv664lUcfw5oVpShJwoSd4qoZA/gVnPnhzPg736TsLmjlr1/tloOWuh4X8iWlxq4bA
XofgExzqmCD7KTTvb7hGTUKgPwnS8+hL3oa7w+O4U/tV/a3dP8gqE+mFDa0kq7lnYFiEokOwcRsD
IFEtNGOsNZxMOJlJbgljVE4xhO+zavlIn5Zy+gkCE3zPAuQ6pUdo6MG58q6RhvjtRAziOVvDkpL8
VEhMDCxVDAN5Ec1j1gCdo9dGY+/AcoAugSHpxi9CUJ36aES+g38dsvyPhkkOBUfSFiVHPsSjR4we
P76dXslMic/eKxb32lHURZYh8svUIU4zUWbiBuvNyH8VRnv6gyB7matAc4kPHqMMoAepyCsy2Q/l
S5BYcuND/+Mr7B2wGzTqd/kTMGHV8bFXnwP+cR5JhC2hBYIvoLby/vkYGkNpbO+b+8SdXAFiKL3j
9HedraHx7Nf9AmQiynCKQtw0Qxb/en3UksxAg4ox5DBCne83mscULoAap7XfuQYjngvsRzFw9lZz
EGiLcPaorXjtkD8FMItk7fgalPWDQeZh9f4ShkEp0lVGbf6w0dNjb1f1meuT0meWaURuRXLfbt8W
EwhPqwo05tZdyT/9v6qSL4RBcnzj/LECWqRixmNvmgR50865fJ+XBD3aC+iWJaaNTxQ/JhOWBM41
Hdn724negwe55S2wXTB55SYNfXdTdBJ0V3TdH08L7o8AydUMPKvvyH85gLT7zmCK+1xIgxIiZea9
7sVd17qN37u/f+LKy9hBqdp0rt9qzZRBodcN+8mORc7+N/8uqlxaLHjp9UMuO2R0iurH7cgP+6/D
T62x3tPGe1hNDv16Q0A/hKurHsV7QfRDodkK3XFY4Z/erW+Nhc7oorH5Ck3SAuRhL+zhucl5SPqn
vz5E3eG+9OLWXaT6PZjCZPtRBkcWgY4tK+r6uoNAd9rLoSlQD6ZY5k9ozd+4P7hrkFF7HlsUpSGD
O3LnurjuVJoarvGkDQNJ6HIPq0X+V7Q3wponrz1PWyOguLuFFiCUaDoXEFYgGCiepy6O5je5Dm+t
3/hTdJVL15GsYLexHy3YwgGpuJVXSlyzBIJIO6cOwUQ7Hsgw6U5iMEBzwep1i9T4VxhNnzeOPWW4
t2GCAYjdb+rUcLL4muArpP8Z7Ec+zkvaPo/QqNNp6Mr0vibipBzYvAaKyh0jR0pjQsnuUY7fYdDV
0jD6lgpMZeSETfqcCxCXyb4zhHrgJ/W+yRmPlAKx3IFA4g7/bZEjXUoX9pxManbN1smxfGgKJqGr
0xaqYu4xfA0J9Or6af25/Ac8yNFDrufAEEg+lFyY0a8ItpV8hia2KqVSm1D0/PgH7yBxjiA5t5vq
394csLt9b8Pjyvnnk1cXrtxj/J9PmhiTPqhYdGdresXU9QxwsokOo9EfPQ0L7su+BeOk48VSBTP1
pP5FRTWRu7Xo9zGtzKLYd+tV/66f57EHBk8WNvdWczBMD++HWPGQ/JHiHuHJfgU+z1B3nVJaZPJR
cjGog7R7q6z1ZtB15fPFdBqJlnuhJpG7YqtvxOn+cgBvNhclX1UpIWo1wdAs6x/LMamqV8O+u0lh
0x4QWu69ouCWe4QUdh9kc9uRYcQoo9E6MgqGTspdRI8yPfGEhpReAkNu3iuMoXBFcCrNZs3M5kLx
KTGtoCwpF2SBc8v1cYCYqYTAoXs0ss818oWCeBBBIXmB9CHJj8wHfgxXUEKN3iQ5c9Xghz7KP2ij
yDkZFhKi2/1jAjLbHRvvGIAk5gasnZeCwGeukw4orLC8hWrUes6gWt2SQngiArl2z48LOxmAYQy0
5y/aTDFsnelv7ock2w7mvyJ8gBoqYJD5vIQEnyLLFBOP/9poEbYpS8akG0G4+VCJavEe28+0UWOZ
i4degXEBiC1FjqZ3hX9K0hxdzgD8U2K03pdEUYW2BkdjNzgmCjoh4+JHPLTMInyDBtVGhrrxuo/S
iypWXbrPCEmEQGuKQZrzMZLDO9zCK1bn65h7zZor5wXvHo7LTVRBLcb3azjab4Wg1saQ4ffzyU1W
zqHAcrrTl7Wxncx/90Q35eroo5By4EEjI8e/wLOuLolglM0bN3zKhW5Rc8Y8pth8qOt90JhPch4X
RvYOSVRiEyyESDGMOBS3iUTeFTn+eQOYVC/l218Ma61aJxHzRfCY8Ql8xQec+oDc4OLz2NEsJ28T
tiTIAYdPc4Iv8fFMzi1sa02Drt8R7jvqWxCSx3L4mkYDIUlj3BNfM69SlUWBJYhfVu+msspcjQlM
Zw8CHJsnCeqK2R2HsyE6b+23r0lHP81sYHhSoHPNIslyqmGPQwaGoPu5rm+TiVv5cXnF2ScPV1wm
j8GJZoIGpKIB5DqFQlMEfOBh5xZCSVgO9bL2yZdzmnZ6h3dxuor8dmGbm8Zk14ZnlwsgjMvZYh5L
RA4MLSdqKjl6/n78dh1s/5bY4M35gkThlDA2/hHeJsKFJGyL+wMuNREUJZrjqL8FoAmxKy58HXA+
X/a6Pu8xoe/Nl+6WpySnb6cJOK8yPaUDn4ioK2njjDDglIHe/EsNGV982cyZtoThISqy2tpDofP+
x3+dblvtKwp0nBsP4OXpE1IeOw2m17eV6iRZaWAP8aabHVMo4b3ccijoB3QTxYRdN3udiqGBymo6
yb3AZzh9NDYEVADaiZYEUzvwCbaVvlm2ddhZv+AmuPFJVw4UNUhSm+cH+SeGeWGhKoIzRL7ENrTZ
fxugcWKGTj6wdhGQNDnEebXhkosxibBAgM3YcJjqQqk8IXA+Dyji0auwC4VHV7FwY6+pAxkJ0b2U
OxgwpXsu97bpDB/VYea5hniepsq4ko5mjmjAlLCTNdlu63npbjXl41JF7iaatLan+fWk1lazJREX
m45P4qIbrcusoQ7QNx+y2Gm1k6FOd2YYb+s3cW8R2foCbTqSOuKbS3HqcTxTSOwu+5iDA+uWLc0c
HwklB/422ebket5q0IJBoxnaHUDAw2yMtou5KZbkhOgFIrNzmv4kHciQUqPlgCnco3fpSn3thVKb
R/jl4s01MetN6+aYh6NFjhZC+R2UjkiyUIjkXo1E35NEdKtMDBlR6N2t/+KDDjgS810vwXEhA1fy
ZrtdA93vFJNIq7FYcrDtwxvG18dZDVFhiucxm479SDjyAvxFELizitYcPxw85dsQ7Npv4m310q4V
YueRCUelmd+HCLVmGy9qkzh5Oe1lFMni23MJjgyqd4Dh7J6rQCtWGk2xyBD7d5cypDIX6KgHBNoS
iYRBK+kgv581T6tmdRIZSJ0fmHoGd3fbFfuvpZv8HK9/SpOW9Da7t+QJLi3LDvCOq+cB8yDQyDGP
Qx5esXpo/rpoU22kEJzpsdq4g/99FkyTuxAp8IJibo/GgLnRS5cNMcRZx91en8egeGxPk+xpelbS
F7yKkRgbzGKnWxsf5NKASm4MY90d4JzWEl+u7hGZhogbEN+JCvV/8zgPrNhrwlK2NvuR/BahZaBu
dTC0hhee+PC7E+l0s9hkK8VeJJl9yb9O+Y7FBlWZZaHV12rAZAEBoLioJImW3zTDuix+qffJfk0e
IjaqCm3QEble9dOLJZ/Os3SlHzKb1qVyMAlZg8xam9T/gZORZWi7hBCLuOksYhez6E7HespFnf4/
SvEupjTn1JIAySYuAK0RKOQEMXGSlZyjhNRzgS3zJArIhyYXjOe5c1oj/RboGDD7OChIohfBfq/D
CcAF+zMGmlVmAxMGElT2fNJzAAtZTuLCuLpPAMXE+IIu9t4yAbSVLxU7rqh4ITQarMMIJJT7lkvw
Lh8wmWkIL0JZXIfFhwLYzZcxvYs+x1NKt/LsXXj42yApe3nY2rMP1WQ3xhMLr2Vt7xmsP+YwNYUy
j7St4RUcMCfxUrdE7HWbZpQyiydFMpxKvCV34SpEigUOh6citTgNXjIDZTRiM0gILvDK/aHr4HqF
e/2uKqn8MBET7HxUPQH0pZ3yVZkBMqrvOUl6Wp12KbKG96MpI9S9GVjfSCKDd1kFBnIWtBWb0WV7
+LsOUeseNrK2aWmYxGYWjtEZBrhGjb23it1Iaug0rVhDg9cE4cc6Jl5sS+Ye8P8ziN9eOk9SbLnx
a7HZZzaoF6Zwt14PgnbBWBayh1sq2yT+MAL4fuBGvTSURceliE/ZM/iTlkKg7pLHWkx8ZLpfPXOa
tpDw3LCwgkDGQa1kGLWOn0i2dfBVuoEXHEyYOkw5Os6OCZmgYFBZeyZtu0XE6OSEeg/7YAgsG7GW
olgeKj+PmGSLRelceJQ48aBfuEwgipCqJkp9I8H02vGUTYzTVHc9Y3P+6yRIM63enPzvjoZlpcqc
SZaM9yFvqXy4kUAKkF2+FR0PeAHt8FrEMTkvJ2nQ/NvEw6Fl+fpkv9ibyzCPK1AFgPJ2I0kZMOJs
YPYuewu5OQqXMuFQ0p0eY1t10tD7PO2KsHlw1T1KxFPZeCsFxTAqc8OVHMpfVNXAwL4uez/aQju1
Xv6HLjLulBRjzGUk00wCQ5c1kH3Mp8AFFYkc8MsTMFgR4M9RSTAkBWnLDeZCNOc8dhk83hDVbP7u
cyjKsXFYqZ9KigowTO2f/pCnvfQoa/6uWXRMsZvA45BCDZMH5LdoFaadPq1K69n614ETidFy4W2o
eXZvo34WqKmx60xkCK4HTGRVjSFh2+p00KVOtVtJqHhfLEJRS+fZjZ+HKZ/HycdHjHsSrHnvb0Sf
JHmhAqW1QJRwjvRsvJwf/7kf5Ie55sBCqdkDv0uK5CXbXrc/hjhGgzEm6MGkDgGdtkKJa+xJUg59
pjYl+lVlfO2BwrkqUZ5M6SGayELqwl2zAwiNoFFv/7detrzyMdXrMDCssjcKUExgdxOxGsrBhEef
Xq4D31nQEHdX1O9K/JoDjhpe8O27sxyJIqvsaZKQT+kIaNSIK4rnFWG4H+SePRluXDTNcmDcghTd
E6no7iMkZH/OLuUZvB+NM/a998YYXdOj+bHtlUfgnA8WaA+RrsSAejmBPdqCOvCau/3E8RFzjPsQ
csd4xgRwzwxNvOBlhg1yHUSDYRE3vJqXOOklnGotdz4K3anwzzgbSMQVp/2wrafk8RJa+Nix/B02
4/ERIyyAXUT5fxtPbAFyj3C8jUjiyOON7VapNMcCyuSmlahSUIYgCYgRYLOaCyRb/0RuHjVybz3u
Rqk/uYZqceLp/7a/Icb3dGCkNLBlooZv1e069A9vt/5PLa9818JQj28IEtyBcphxXqd8lIn7o9tt
0IqQF3/I8VDkL//dW3Np5/og6betW+z58Xy/qOo1SWEop1Gw4tWLbHU0daSAOCkx/Qwbfd8fW6AR
+vB233EdbDTO6wcmGzGALuna5jBGHU82tw0FaMrCB1WQqaTlszeVCfuAYAFCsq33MNUtIKY69erD
VkV+DfJLNE6XZropH3ySLRQOqKZoZn59+VLqT+XEvFtTzx5vzAs0dr+mKMnRbS+YJea8Xj5vwmK5
Bo7Gk6460Z76XsfULKfYFRaua61bFHKNtcqBq4MyP3pgisyLwo6tbvKK3lYsXd7bSiD+ZQFVvN3U
rxGHH7vyvfzIA8LqmJ5Nb/83HDb575gEAxGf+bQh/3OMyeq8V1g9xiChGm8rHO4sRd2CqKZn5x6A
54VZwsdL2UvzkboRSFp30FaNxh5bg0yTA0ZaumKZXBHyNMvQCorReaXbYAYJCYyHXTmnp87yEreP
x2H8WMS8ygRA4QA46WMw3NPONxVLryHF7sJb9KICwXZGQz0LqQxJDG3+ddDtNKSOebTDDrIt2KoS
qNJsNM2NvcBlMQbT29/+Ga+8CALHkAcnojpYg2aaSe7F512TlPx87H80isdZ78vScJCuNWIWgXlQ
Iur1I0Ny4P/kEEIBfOKVuejoXgZBRtngZ6EGE+nKa1e09BhgdfNCJtlS2P2rzhxy4fkklf6MYBMU
JrrbFWNxjoCLZD9UDORXTzsUTdHRMToCgLLq1VoJwmbXrRm3POTQRoW4VuKViGd7J2cfTqE2g4me
acovAK8P9IXLTzdKWNE98fd3FBkCvoF3ZS/2zwZx4/ckpjDssw83d3MK85nOyErq1WBy/gHjr+gf
6545C5fzmNuQ5HEDkvLUGJpIH+qHBP6eFmgd0zjJk8TXqKRQqGLa8EREkNJ9mS2OWtZHaaNHionq
zczxDsumTAY+CIzqQdfRDHXepjfLM0DzWU/48D2ixRIZnEnSZZSmW0DZTfCxfsXQmSbtRDcO6hzJ
J7159z9jREoPYR17Ko2/tm+b66ai9rKq77j+FBhVUPn3OprFzAEIVDg2VAArl7xnyxKDDXzaxKwT
9tNvKrdos5LEEyLPAlhNexbTUKfKljK1GahgGiuAWz/8w48gD29kf9K50X1EHi0pGVuxJ6y+srbg
P1zbpquvKuYYf6Pg5qVj8KNY8zh1MqsAOg0zlgza4GFR2Psdrot6B9j/DXedp+ieFxIjJ8N65dH0
gu/Zivcr4lDFU2tC3BJtGDE7QBd2RQ2UMPCkxWnRTx/R9cxf8xpKVl5GHoBb7a5gQ7zfqLiioQWB
ab9WFlaylprWb9pJufL/gf2dABwhYlgamdIyEz0Hu6f3LuAkt07/3ZutISHmUM4ki03TCmqtFxUe
tAmmQ8bcS6UVGQhLRcBZ5yMr+lRV+U1FjGb5J14kg5EG2J5YSvyY1c+MHznN9LyObvgVWvvn3XcG
QxW6NReyAikURj/9jQsHO21WstdnosQzmFtkxNceJGlxtC0Gbabrqles1CxGIvMDgZVmV4goweij
L3X64jNPw5oqQ1/xiB1ALkL7FoREKZLHtCM3wbRryK/+BKedZQZONC5j+hp11zrrHpiXk94QfS4a
nZAQXr66twRsxMYx+oriVtUUyiGB4w39YvKWLfefnPhG+ShkMKaHHShMNUALkY48K1XuWdQTvqdD
MCdHxgwwyiYIGunAU8TsAQjsQusjLlAFKRWlJsTyJ5OtFzEjE6GrwLnnnp91b6sNLCv3by8PrOBo
SXbEV1O9LBsyEcw3M94LYmAozu2vUWWpd9ICltqPECOFyEAtUjxEe5U0ZczM+MoCx8kNzazJVqIT
NKmcttcxKibRq4iwlm10vNJk0ipBytH2GrH6wGqR/UFH9cBUfT3uCRTtZM4fZFvKAI4LDOdV3M+K
YA3KUkihWq+XcQLep4wyO4fZUFu9wuh9KielAoDzZm8/LDaDMO8fh/SSjzlKVXkU3D5nArV8gEII
P8qxvxzsr2qXpfVgZi391bq7p9vpuM29HJ9pFWNk/qswNQ171jEE69UkuCf7YJKR3xMV9x1AENc1
e7rDASBBUpEEpomVd3+YU5gbimjPfAhMia5Odh0/mkeJTR2KQhUrRkB1jmrWdkhjxzr60r9TeIf+
6XKEq9UadUkNA6sfE6KMdEbkS4J+6ZVwyfJFb14QUVQxaEuHIT/hnV5C5mHOCdY/6OscCAXtrnMh
FAc+5NeTIVfOLUSIDnUBt90u48OGCIYbiHUVu/I+ou96/m3LbWsarduA54Oc4CIymyde31dHsRAv
jikj7VMhhBbE6W4Yow/N32KOgTTt+25sP7/X1olCt+c8hroZMraJxXFqS29Enj6bSxke7gfkz2jB
arlgkIKQPlsuEKSbKpDU7ApY48dwoJvIVnBwL8/JdUw5/w3X6Ipty5ottkjzLIWm+RusseMigShn
An3btBn1Eg8XtxPk2AfDkix9a1UMf3W7AgOGYyyxOXddkueidRI3cTzh7WdQgd6dS8t7vCBYWCDP
5LwUge983rnDeynUW+iXzFSQI6rjY9rdpHZ83FGZFBD54QCOYIxzwxv5oxJF4U/pCl1ObypXQ/YP
d9Ed75GsUgJblTKZBnc43GEl1vTvlTtHlSpRqB5sVxoGtokATcCQs1W9C7SwJOQZYR00NLmA5UNM
kWXATrZwDFtNhdi1No9soxqBqlO3tfZj97x1JldI4mwGy9dmTlGzNLRAfQxEysht8b5rfm+rHMCn
H373EPudmpFSZm1fI4S2PaR0bPF5tDR6l/Z23SIXklcZQRsgZ0/f4kWunCjEzwc9ERKA37EDU7f5
9n2Dar1rPAbvybtDBQy7RnIVWCtv0KZkq+sJVeXLIlRZVuPFZB7ijXOeG0LSaiHcsk1kB/F3EFNe
iaGCM2KjRLB8kF+2TNGUyD2wPbBxfcwv6z2BWIG6QXLM1+UAFaYaZiVAMnwuiXEnL+XWK7SfrzTi
cfOj4qK7VvtUhu4eSIQ4mpTtc+kaOapSg15AkGVjaA/SOVBIYBoT1VG1CJ0Ddy2u8MqFEtcx+pAL
8wIYQA8k5KjSV50R8jrAf6nFecm/nF92g6Uq5Wz8rktNlny4hUuvYnCaRcOp4U7GeFXWzybl6+AS
WkprGPvfB7F4ob3WPXAKrqAXely0dP62QEl5YlnbUR0OE+XnMUcJhLVbpgPW0qJrkDF4iu9avQDT
tAy+PBo7TmxsCawBB43ysv1U8ncFDMGAmu/ChLD7pe5MvwKgJEVhJ+5NU2FW44KAMvl5aWQp7ziK
FV6DnufgcT40CmoZGpZfp4K22NHAd0tnTh7I8Dqe6C6oOtcrutPOZjzqAh8h5SYos3hMEMHZgmIN
qGtm47aZgYGDNbSUWEWGxtorHGCHIICx7fknygwhmqKiCkGoj8kwQQucvIHbLx5pRK/k7LJLr6d7
HIwS7B8Sgpwu6lO5jN7AxXYtgFxLQsyRbeHTaYS6j85rGkB+qgSGYqEB/ukVo9rlIOAGJHHJnolj
MCVkuNOVwc9SwSRwLqqbuB3Dp2xHs1VhSWnnenC5wdfWyj33V/i+ao5IC/BaBJJH46m+evOf3Rb9
Sm9vxznmuHW80A8cq/qPwuYLo28ImITnh5hB8SdLHISFI6GqNqpv3Qv1+t+NvrWTOsYtH478QGPw
6CQ4K20679mWrG3r8ln1/tHlHmu/4HIrnBiczsXOhqwJTtFjjrhl5863wErSLjzkmrfzQElKzgZe
41xkMj4gVqESHE0LALVKT+ox5LeQNZXj3liXeLRXvVZ0WzOpiVq38B+yVXhpCbZotmu0844sVllv
ZrnnWCNZJNyNicHzvYJ4nRZP9eN3pZuMt/QJjufdLaJHs1Z+RDU3S42gzbr4cJlWjLeRsI6rRYM3
CXBcfWDuQ/Kr+9X+kuVgL9pyP2PPoLm7ICidmaVz7hML+PZ8hoF9T19eEPRQayGxpRp8ZL7iNewU
zQwwOTWLBJ/16QlMRZVi880TT9nXOUZqhONV3ZTRp3ifO4/zIBtEcVyZxqmUYCFUodlywBI1JzHo
VqnJXfRbFRMOxBD46PZoOZnJygs64hCzhsIbEeuYdM68DG5hZffDUDEYQqo92MudSOBcmxaAmNsG
07Y6o+po0bb9KLxK9p75ldk0qdr1A+UlZXhWiiphj0HdKJ1+9DrTYd1WLFoj2p2S4HdYPyUR795w
ZRHoiR0NCf9PX24pLslRTDNWDva/15jWk4E5wTPe15at5qgBfNry/+TmeeAzhx6q9xN3Z0EAuWC+
F7JOgZRuTUXGmYknmvdedMojsJEACuahtJiAz8nPrWaH96if1UgnmG7j0KIHuWPFLtEE9UWfTdi9
WRnhN3SyFyx5j29ZbMajSxg+3Q6fG0k+CqBzjjVATtkC/2GyU5JyFRXRtZHNhtuU5+dnxQAX6vk6
yiiC+Yfg5kVuG3q7puwAYfRZEVCnfU8bQpijQr+03gFkLJGke6+LMCPORmzbkBoi/riSs//Pzitf
TonVxYiOtMyLwvVNRo7FWxGUa3ql8HDmDxo8ijl5Pt0KzJVUlekI0a76UojQGebuHir1r5Npun7T
Mpfzewl/FXuVNOYGWfurEa3li6T2/XHXcIVmhpSk9gAlqE+mczM6S8VAmhtZA41TR1mHV/hLuGok
TghBLlNOejWyFPCkQ5omp7R0s1PjfJ6+UQ+aWoFuk3Ii/ePADiJsyizSSaLhpFtA7GE+ItyuLyhg
0s1kZ722gbZ5BRJzShQGRiB9b7gW8ntCe4WBj3YiKKwLXSVoXJOyhErunCSmDPOhrJVO0LfxDlW5
w589pnHuOc43iMGVOs2w4WombcbcwmFvIjzcaQqTFIJSUNpKGk1SHwD6Ea48OcrV84dC5D4XbyfE
0ug+KfzC3gnMA8DZLKuHB1pAYCgOhhs3xUsD3f9pY2mkzXufTJuxngMat5PesVMvkSuxcflzvYb/
a9FxQF/LKdQ26lil8U7JbOo6n2C8mpCZmlc5oZwTqGCUfvUe96jHGNIytOJORbADnak/UrkKi0IZ
I61isEoOCZrsCHl8gb6JBHntnj79ZmFGrGrCohzaMmCAUvDjW5Dur3l1gEi9VzfekeeXaGt+fT0q
K2Zp7jJqVkDkHvAm8WykajpOUKE2HxAaCNWJvB/y2yPFogxCp/brHIwmoRKljIgX+OSEJmaL07fc
tqCk4uFOp+JcJr1HQ9k1a58fwGpw6spzCvMHeVIOQ4GsngiC+wmDuoh2hrsiLHZASfsKMgZNdh39
kxUMts1z8cqAhDhIDqO5e+OTDFdMlM4lMKP6sYv5GmZ5q0FZ9cfUWN2NunlZhPpCqVakbyi6apQS
vbqwa9XZs31OzRH07dFYBMTaSBClxl2fkES1PcXXgcY+mLWcmkOb+X2FR98zPaytLZcEia4m+9ml
Mn/lFGUQApFbHO658h+5odIxPG626/YT2ro5jO6TZTTdUebOk3KO3yuuCEOCGsxV5uKarlC36KBj
sfhb5pFttVUsh1Yo351smymQjKJ91c01ojI7Zq4BSz/nCVsWLzwXyYVvH7lr+wUksFal9Y2YX1VG
OxQlNQaiRNHls6naX8BMjZbUIYX6xeTIkgYhUv0aw0gXuQHzSMg5jgaO3/QbtzXtf/38CER39zZ/
pgDSGVoxCLk6Ps03jbG5Znz24VY6ddUxCN7Ta7YtrBKbx9WnKeicGbsZO3sQNsdTKYEKIlF3r1fu
jBwwwgxrT60byry0Xe+uClGFUU5Cpa9e2uHusfuK+HpuYWer6jRaI0Pv024L+nU05mA6By2rILgS
C7SihuGce+DMu69TrY3RB1kT+TRqkX4aGMBfwE7J49uMY0KFS+IVQgPn1GydnFlKGRWI3toavkHN
Qkv0fLPVeS3rRuW8qpOhnMqQvrUDkRKwutO4bQygSuOPkyNk698i2+1Koy2pLG4Yf0SpIhAVcOl8
+SnfxB1q9xAM+MDc9UXn2ATRBvvlDpYY8strUrMQmpfj6Z7e/7y9oMuERVv4XpLzhThJFWyNDZZU
UFd1mVsuqew2jdP0JXbxxxri2FgHA/uJ+HY6ucG6BkM7Wn2JgF5SGAme0x92yP4KOCobuG4Zo4jN
mPQzmyyKVFf1cK1ybMe1gSyVQQj2SF4AHGXxyR+ckkFRLeTIq0EeXox1kg+0NewXIzI+F2zycoxR
w5si7hAd0wQl9Jb0IARWBEYaQLIXH2oF1okoB+Ptj4EXJqYnr8PvTXKvAEfSdYo3WBL3dEydk1Xu
Iymp95B8xIkujNcOlYkLNR9ULCo44idB4qzBZLyAkAksNwrt/P756ymARsVczW/BOmDNJ/8CcDqR
JcZqJHFpv/LeQSPtYACQI5TaWUC7LJlEFqergT8kqbqulVMfFx9qpGWpew9raqSKvoIDi+fpi/7O
R8FX4nVJfa7OrwFFz5qrH+eR0h0/ZA0xzHQEqZoizc4gegyX2d7w4cmZeiT31P5x9qIpGGCnEiES
kraMV7sCsEtfeKbUU0vgWsHeNl4HXA/5ZVPZGxe01EIDB7kyRlVWAb4eNtl/NsyvHxDdDLmXBFlk
4+EqlwB+XyBbwHLEN81wRt4EbisnFGXsbNNO2/kK0oIk2BBp0IsI9U+Q55hIzikagzsy4i4XQ4/v
64qRynqH8/tQ+1q1EKCrYEx/wM0mK99qzw2FFjRT+amf3xI/ONUzAA1fXJVGsVNFrs6f1rpbJEll
zxEKcHXaQ5FUpX2umsdf+RKFyD5vhRjMHigwmk/bnmgdI9/vdLX0tHFzyN5TRuZaMnTGVzCO04qE
Sfa09y4vwLpdzf9Ijp89MfLXrLG6dl3zX+0JJdtQwGvoaT9N2qi1gGuD530D6WAwKPneeKpjmTZ7
Ie3HN48qrDiH/tjaiB3E+U1VOK/i6EhavLVrPMy9DhiY9iSS/UiAWAsAIrhQMxL7FDPQkRILeZEN
HW6l8kc1DhRCEH78K+rWMGh1dX+ZeNzFXAD9QyUBQRelDbeIbCneoqPTZ+3TFv4DYmDh9f2um6QG
rTIfDNQTFDd4AfOJCrHmEjMFCoa2SHeYCdLzg3fdoeLetXjHE0VVF0vfIv8l64F3R365erhhANCF
rlio/EttYsnsEYKZX+zcimZ3x+zpNGm0MPwwNyk6JuNW50293LBBsKmYpMhaBLusyNLGRyyoQ+PA
1LqNxrLY2TTOFifpTVahnO04HuNgjerW7vs0Bkf7ZzQTceE7lCeD+uDtchSnllTsH3O8bKUT9eqx
VnVFblBp/7sHrub9jTStHWctluw/MSTneYZGIecgc2Y/F3h6FPs9MNw1iXYUUZk1G5LqGPucthHA
8ThX/JK2SjlTXa2ju9rcth7swnBCAYbX5YhG9pyHMomKfmh08Jmxz5q95uaFrcVNRmoHH6pTdu+/
f7G48y+Kh9dFuMBFHdHNs9KTOYooqIeFECVP7fV6mePeX88hpeQK0dVu2E8c+rP3CcQZq3w5CyZk
jzLYmTYC1g5IbB068JqLEQ==
`pragma protect end_protected
