// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
ZH/y6qKa+vlrllRWPznh0Dw6i9HBhi2Y8eLL1BXWxG7vGZpe/ERv06D/Mgzp4/rFYxt+N5wrNrhD
2MM24Vg+5YX8se9tbsu9R3vxU0NfS7RKpc8Vk97NqEY4OZ5asUQJwHrbMoBuRXK1HxNs/ay1w/1W
jEuOqVMut8PNVThhHvKbHRF/KNlp5cGrb7YDIKCwqSqwCB7Yv5L7yZrni7J+U4kDDaxaN2oa5XAN
06a3I0EYS1hdfnkwUoRIl+mHEAPTIKcBeFtLsj8fTpZ4H56wiAhPdcMRkB+MrZHX/PAiJAv11Fpd
bCPKtHhwhoGSTL0ly8RVzAwZGmKbvnlkcLJXwA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
IupVpgr6CvhnCWrhCl+LQ5ZbzPapCOnmjN54SGZ7e3ZpiXgCjyUGus4IntCeOOgMuMJWikpKKea2
ljEfcpFxpcHic71W/QfoBuPDNQH1z6vJ8RdwrcccvLBhrPfuxV0SzEOBofdisSE2Ydw4iUgkhclg
hqcPUAbqkz5/4PDKga+v4IkM+sNIqtG3Ey117KQHMr3zsohum8Qa5oq+nekos9FsHzB06o7ligWM
uGpW82mtCNihk1mLExbecl2t1kPFINweAqioffQsmDwlgyac0evbrIT/iO0lSmAA8Xi4yIyR9PYH
t9U/adDo182YkNI5NuL8MPjazxouNoplcgtmNR1lJ6t+qZ5/cyL2+tt4FOV1n5/PVp8SA60xOeSt
V8XoNPQvG5y/2zhaUYJ+kLoIE5aI802QlwIQVVvDmib/013xsP+TFrLUwykwsTDbZQE5Tx/wd2Cx
oXloSFWSKDnnJA77Tw8wDrdICLpDkY/oIkIDhNT8itqMzSbaWxK+1TJUzjsl0UUyGrSYdF/Jxdtf
G2HL/lb3a1RpXR5xTMAoiOI25JZZptGCtIXrGRdtAJSYkT3V4eE8i+/CStU8UULffDq0+vXNm66R
tn6sYXYFc7XqJbRbfKY8iVqKwcf7aVMOC8MfXWqvSVdZDMPd3UnycGyV8+BiEOHZqltsQjgGMPRt
+DyOqqG0PxFXs1/8ScWa0XNBKBFjecpjzH0G2sH+wvITAeCim3xxPW+P8oeDVdIO0G03cVf7OB1N
LL2UIa4mDoPwlmQVRvZ7ResT5VJ5GthJPf4q8TMIWrRPOeuw3nl70PojVnL1izxwPNq5EIou13Hm
rEGEByx2KZl9e7aOKQX6HGUPTD+bUfJ1c8Q7TOtJtrVYJPRkmc3/3nFGR8VvM0qMkacnflP9U++b
GVbVRI7jSwhrb+RO/oStDMbcI/5SFnr7XrkmcJ7a0NhF4TQjqKbMxfKAVRdpOI1ZZ9qFwyYV8WG/
ATM1Jy2bCwEaI9qRCypWu559Wbf+6odvdBX91Ea9sAolmoi6kswlTVhvHxqhAmCEbLPM4k7pDJb4
wKJLk3ll7dqsRwe8VVNo3uj2zzgUUSvpWEnsGBdPkhkENRnAKW5TWNlPlc9N8jhHZLQV7lcfcl9i
qcnx/gYF1wnKZbZbBTNkrBeWsj6PsscwYruF3DfDDXTnYswzPBhTNEs4AQhB35wGFxmk5Sbgngnm
nyZMB53e/nNsM45LSCLCqjFgjKcFMQvIatlx7hnaWO8iEqAqNfrZ6Dv8Txuad1pqyjBUnsdKTqgt
YaVG2ismRjyUGcBn9aTHu1kBNOze1NrezfoPJrLSiDwSI9GRJxkbNGZnVJrhMdLWROCxvmAhzzxi
iBSixLauvA1mjJk6jeXLlzzbGlQUkSx6PVmFkAhMByLAd4haacjoZavwYH4eAiyzfwvPiCzXWPug
pTBMQPmdvHuU/7jFMkHSsrEJ2ui//S3CXgg/ONOqGYZJ1a4NvVJNuf7UXoBAh9guR4sMtqv9oNi2
0zKIPQJpu7TCoikaqh0PBq4kV91grOJp0GlnqykrfalyxqprDXe5c7Rq9gJ0li4tsh0h0X9UuJWz
Lj33N07uBXaKfNDuCejKktojTuqxR8ctCVOg37uEQDTj6JJFLevRIm4WQxOmK2fHlleOEr3rH71D
TQjUnXxiuIZ0j0vG/Oc1IOGDRUFgrwLmDl2AY6tPc4xEvgLCmPcxVwZh9+9dCWydXheVcX/aEqD9
4xvA7BkvVbqXoulbgOfMcJZIa1YA5Fqt8oAlPEGvxjck6QD52uto34Vn7k5DU5m/Gst3rZ6sBCQa
2yscAF/YS87Ujn4y/yIiuncUv4OozM/36tDMFV6kzl7ZOs7YDHvixi4WiBQUP5WMli8U8K3SoxfW
Ng9WgyieHwck18nhIy5VClcwIwb1d0OzNEa5+AjO/sy7O4d+qXVZAOnM2Cwrk5Wh16ZkmaDSszlk
buxB0IEKJwVAKMphC3OWpPpfX+xVzTIm30IVSiwUUQvrCXXUfNVVzUeceFXZsRXXAOcDenEJ7T11
xWcwkTFmPxjfqPNlerHWENEKow2dXnlsRjIkQVzuRLtUm+v51Y0SXsYGa0i2LHjgBGNhS2RjuFvc
j8XuKKu3OI1S9H/yd64XmKVjMQ6U/My+RTnFEg6U3IXUIBcpB+w2CxHAFytRtuM6DFeGob4m+n53
B3NKNxwg4ts8UYsp+30EQfX+d3dG1L9jisGVx3vruRFconqn7k5y9cONw91iQCpTWSQeCgVibths
ugVFLj0cDaImS+f05wrOO1HQwNqtx3jl0zHmCyVFBmf160y64G3dfkPLCEJ3GS+jG2pM21koWjtS
VL0QCUUp8iGsQhUW+PgdVJraKRUnk4Ez2O++9x0MN01L2jEn8JZjM6dDyW3dnjJPZxTu565A3go8
9fRtyJM2ANduXepjygh/wFKg1ojdXLO9airfwF4eYS8lKH6nEe2NJROO3fu/S7VeoR5I4dXqgdgG
xfk4NuHAYk/RZmWf4u5BrcpqS31C98RYR140pLJDf0HsXhpKd1CLjxMM5+LcXk3KtLv44rBKlt2+
wmeIK6Gw4vNSXgq96kKz0a4Y72m+8oba4tULumfqUOKrGxSH9h+qO57CaaUMnW7/M1ThAC7+nE0x
/nJwtOi0+F2rkU4E60Qhcis+8KtzYOB+Xf3ptEB6zorH+8owVsqomu6fmn1bY/hnPO6gQeIRHTZw
t+lxzVSjLzyJrv0NQTaG3PFkcBlhpr1R4ITNi/t9YMb6zAAZP/863vKiRhuMY+KK7WLhgFfJYhu3
sb1fXFqKzLlv9AUMBVv30xp7I7rLmKK5vSilgq81RH/Mt5W5z+LFA64aDPAUt+jUhu476doWqzHy
zVLAhkdKj/ZQeEM0xGQiDWBqE6XPYoXee2HpX3BZuLJlTmyR2bTkY7I3VFiSnoeCzrvWDWOXypmy
bObQDQ68ixr2McZ5w+Yx5XrZDLMDoctyQadD+kpOTNf+fjh5LeQESxAQe2DMH+E5BRP8rnRDCXX8
kgBbQ0C3XFpcH+Wm/y8iYVzg/ORKFSHiP7r09aK61LwupzvssoB7tQASWtPYl2uoa8Bj8jm6Mto/
0ewHxcZwTN2m2U04p0hbO0PVT0oyN/4JC2IDZ/tGrv9Do/nBfhEqLDhQXPKLlz6Jpey5UfrAgxm7
AW/sJAKpyaafen2VbDWpkPFTQYIuM5/cxRrmfRJSkTjpQQpBRrOv1sGhGgmgg5w4jJwrCEsS9j7b
lIjhx1XNKu2orukBObf2wYarprD1wgtcYVvM0CKblyKNqRh07LgxG1aNdJ66i+djmtyip2EbCj0e
HfXjkwdSOBn5XiXKweRw81sFwfABvjo03VFzO3lfgxvvtEoMNlmynx/qqTcaxV8kNd+3Q4NDE9YC
PCny0XhxJPQufUuHmdlqs4pFl/DjU28iuF+2ye/DI7I+tZNZ7/6idWQQoXmJF4i9u5XFrHLEagE8
8TmNZ6Yfkyq9RPICTx4JfdzFs3424q9g/uCgN3TKjbCc1WrGPEMXjgov92FrS+BXpO1Edq5JxvFq
CO1VPZQ9CxiTkUo1DaxGiWXoYFI5GT8cDs/sVCwBNbZsRN07uemeL8vOeABWlYjEmhgPYzGRlDJO
6AOsP1VCnxJ7h+DpQ6S6nhpyL9NAcrs7sIokgsdTej9Bwt7BxpIcUAsOw4cRYa0jn5k2h3ZM5cA9
TK9ocsDxQFgaQf//7j6/AwKi7xu0+3wxdL4ZBRcXGy87xb28YLe74bh3J8U14/+OsHRE+GhF0rvE
DOTVzkAlkN3u7sgyrdcNjvIvzujPUvZQnXRafv8Ihfb3qz3eSiwLCudYHKkP2/+c4Tfhg0P1r5qZ
WkbBngM2LpCmhQ2fgx5K0q8VxTCSUvbbwWzCbS7seCKhK34HwrnKFQ5zW4w2IUXXDfmMWxGORIdW
MN5i6uKp/+T+6vF933U65gNh8o9bonT3fvReIs+3U7S9ObUs4xKH+FTMH6qJYfF2l8fUTjcv8+xB
dR3a+xW0apA/XlDE7VBIxUye2gbSBiNMwuHUc9VfI7ojY4qYC4SnBXJTfuUWzSiAUCC9kNPhXGW/
h4q6wxgAbAImceSvWHkj0Zq2Bz1iJrxG56BMaMOibUd0Qapw23sMQ2wkahHMC96yvdnO6nMmcjEI
KjewhsPwOjQvugLL2UUQLt8Czg0yUP8ZRBaxaNbMUxTQbXEboX9c6S9Tfb/SHqjXzJ4T5VbbRdqF
QCAmvto+vBgr3BakwB+PCNWnf8Pyl2qpeqQ8+ilqM25l8KYEXjqJAmgc+aT8iS/kq7zIH5AUAy4f
LGElwjUOU/4mG4F9wZH0xwdzy4xfIZpHGIIQaT+OWy0UDmPQ8v4imyahFUZn+gPOcJg7xiULJ+rF
UFnoNm2i7wFY9tkiTYhclXFrea0W0JLbtXetdYFY0sGD67CkKFKM6fY7F6w3VupzaomQVX52wj/G
1C5/2ks7Bg5eaB6iqmuPAmZXIMQrR2XOxJQ0TqBl0uMJUIISF7vm2NFJrCITXtRiHNBInuYTv7Uh
uLJ0JD45yuuujOAVDBOUVeYo6YJeHDLexMGsYmaFLUPnoinPQdHB70GZ6mJJ55yg/Wcg3KbOtjQ1
hZXPMkUaf2qzreN+tChEFYpx+Nsrb8TYXE8zsIzq0x3fbDMkH4NB01pA3mH4MI/YjR90DD7YisKE
Lkb50uJDmwM1QDOqhWuNu5KV+Ap2sk63a2bvVE+t4g5hBhPEvNEtrSOUxwHn6gJHhoONqThfrHVG
zAdCvlEgWrBbqACV/zTMmXka4dA+9E/FMs1kd1scJE5TAGpfQ24FiQPBVqw2oUAsNEKRuQqz5Quu
9DAurhWKoDBpbvOGBnypRaBKZ/jpE3elvmQlTJA7KWzTRKN5+e7Mzwe5/BsNu9Wv5OMZkcSiqU2E
m8rdvUbJ/q1YvH9/LfvSTm2bUI1Eq49PLs0wYbpIVVoWMiY6F2lz9bVgQEL/KRxAV8lxgsezuvnn
wSHwMPWV/RtaVnc7716Ab3Mfj+f6W0Rcakn9Jbh9/VAL5ey1omjVv8531IXu9FYFp1ZeF9N6eRur
EgQc4n0OBatA+uKqxw0WOLa71X6QGn7bd9wSTm7NhchXhlyoIE0SHBARyA9cZc+QhWYXqERdI78I
5PegNJAYpPQWVrM9UrIx4KLQLggViMKBh7hhWvfAuhM4Qs+od6eYq9Y5HwwFP+hLAqNbdHnRkvnh
oom8E9XDekZ7OzbVfg9/D07JlozcmHl5DkvR+ec8MCmH+Av+RvPXTsfSOW4XrNUIKwyje86g65iH
boBqjk5UXsLMamsUKUdzmDqMTEiUBUVvGbTAvSDNn6D2+TxE5ZqJrtOh/gx/9bv7YSwwPHwFOh2B
OtR2lBCNRq3iqDIEdzTZygFmSeYtPRhVz15f/FPeqzHIZX3pQvaUnnwigHQ2VJWq7FO/Emyui/iG
6TJ2afWFycfd7JllopdAeFSeKkl/f0cSal+RaXHZSDUk42BSTsL3SfBrpXGzpr8LDNrB6Eco5R6v
uzbwnPSQvfMy+W2DmRHHcQRYx45P2VU0wAoqVjte6IOZD59oQZFfeu22FUcDlO6vaNmEnUYbsZ70
T7tje3c/XAkdchLS4x4NRoIiQVXHl5wy487mSI2bFLp6bba1HXRXd3FhgKkainXsx7hsTOV37Hi3
fLd2RpI7WvAAoyRi5pSNFojNPL2rNcAu14MRjnqr/izsVN5ozvu4scv1yyzqS7bA1EGr2R1XZtbH
8XFE4gGRonWPTc6F9Z5Zd3MkMMXnVe/xJSI8fWj2FdV6rm8qhIhYYPOmYSrCqQT5AVVQxrbQBA1c
AgOv5DCCIo+zis2LVvC0QdQsBgkXEg7kCfjlc1SQcd/QqGRF2uF2fL/DpiokufN0fSgDRDFxIzKj
0jYfJ4sqIxXw0kCjZ26tTGvEHG3f9Lq2BBVk5+cX7Zj0Sec1gEZlNbRE0Fjthro8ziYjPucIHJLY
pUqBUkLaXCHc3D2CByc/sOToTFnSSP52h7JzjW1pZsjW2jaLl5KXp0rtVn7Rp8JSYDeqq6Q6kpFZ
x/5pE15iqdn6hw3FMEBaUIb7NqkTJZztsM/ICpYKu4ACEbM8dne2WNj46sUTDz/mG5aQhryaxWGW
BaYAVVcZux7jxY3isUB6HbVpNfBK/bJAUhdohEaRIWkixdDV7hvsc9Gev7KbtopztDW50akwwFyb
QjymVtNGouJbeWeH97o62//qVbddTSFI9S/OLvC4yVKxxcQ2TM7aPmzjZjj28tTTFFEJKdXOnIc3
Xj71rO0I1OMMD2CndbSn3CDGwrBXSysDDx5iWBM6aVruV/6ciX+e8AX+EiYuICwR8cgxflsvTTyX
u387fOh1IVD+kAVyshSozTlFXyETjHPtc+sWrEYa+cl57dt/TiKYciVS5BYY2lS7UdlyJFSdPTc1
c4O4eHaLj8G1R+pE9AntFcIau+TzizWsYB9nxXfL03rseC+mCcjXtRxk+oL/rWxmdWr7wNv/sZe3
DSNB+o5HHB2/cAN10t+LaEkp4w0MKb7tTbe5NKdVJz8R8xiolPaKtDDv7XX8w3lloQuIB51fxUC9
zT17qqzcNKVSFXJ4bo0BHCi/XoC40pIWqkK8IBE+hZfMhcPLSe+UdFF7Geo2+KDMaHBUKs+krdXb
bQQYkoZjRlimebktUGIbefbAXg2IlhzYHtivsD+SdDOqE5xAhsBXYMD3SPXyyzuQM6pyIJyAuT1K
9xrWzWcLofKwfM8y5qZVPl1wp++wCnwRceY+FfBrxGjuUVYb6M6UOp4bSwNyX1Uw3AQD6j2NHcPx
nWvlvgADRiOf6HSiDRCkBSdc8jMMbEB9w1gut+F5Ua5I9rtZ1leJXtJ9n4i13NDk6/i1uZpqZ18g
YsOBCTwyYgJiO3ASAXx3gCSyNZeVG7+8Z8iPVKOvA5RZjSyyLIJshPik4A2hwcWw85t0w8kcL38J
40T8nt2w64z3E7o+DV18HOWJIuBJfNgJ+M8ysmcEA8uFfU3nNBQ8OhJgPhXzUX6Wv9v0BAP35TyS
fxcExjfZKLxqCIIQ4FBAAJCuzwDviy4e7LceKv1sPrEBtl6aUQKcH0O2fpfOvDT6j521USTdFxiA
OMZdBElwP1ZlMm1dZUNi2KCainmvLM3tR1ZG381+ElV5kKFEA1+MbMCDT+yHk87a0JBp5WVpmsvb
Eiqo3sTeQtEoOcI21xQWu6I6QYyXLGqQbZszV0qfpoPBSe2N1vN9y1EHD76QrJ8/iJVpCo/+73hn
CvoNeTkdNFWQDFjozEMsE7bxAGrDKxhoJZbSCBMhralD0swy3uSPrfNczgqa/vq+M00EqjhYSioI
kf0ReDyjYQ7z6s+QU6a3uYMD+Yuo2p2Sf/CsD5HRqRLXfz7ds70dv0h/9uA3IZXe5AfRRNZX39ut
yWy0Kmqn457MzEth2PU6gzKJl3CqZVnn41L7W9Ecg8jC8WGyri+e5b3A3VCLEaSHdLGPwdxM3ohC
6DiiiEoIDDo2l/BEYoE4DZtOTDdLyR/kxFJJ8mVUfEnl4gZQDH8kWtiy+zrpjvJnbQ7yce+Z4vU+
HK5u4DyKLElfyv0ZG/4WQCtT9vFWLcBd6aUInnYCxR0eEP3cv7Dc12xPCwL7SMlZoNf6na8sz0a2
Ac8+mnrYqtvuL7Ow46Y+JuJjzc2I/WXL+xyWHWN2LDKW7BAE2HURLF6eLvvMQ4Xnv3tgaEbjjeyv
I/SVq8hUoRrdGnksIrU1GaaIOXE9Fmr6Xva5m+W6ds5Fbk4UrzP+seV5jflvKyTb6mcO2IzxqRYW
//m2WZ7SaUpZ1U94D1y3Ul8aPZUbXwDtstxENFWFokON8FttuowQqlddLwwm4q8135ZdjAEy6Yyb
FqRhW5mUkHvJWYyIZDzOyxLaURG8L1ro6XFg8t8VWWNzWGIC5WTJO6u08MEiPkm1L2GT3qn1y/7d
+fy5cQ5NP5m91R4W3EZbo8kwMKBQYN/s+HFaUoMaCyrIhpOLeLYSZz0qjID7VTw9hc8CNHJbf5L4
PGKm3w2xlNL1fbJuRxlDlDpLZRRnJDCNDXwzwbix8pwUTN3zC0tZHZxhKcFknoAmtX5h3jgx72r9
4voRtTSyrIcIvPZCP4BUA7/okkzxDpr2LC3tYVY7rJabDoXYmTtRYBjpXqcmz5mKzLQ2n4rhsJA5
JUSZnSCK3xWu+eHBYZ5BvJGI60Puy99RVUtxR8urr52x7ro3mbfP1l6Yk/KA9Y5EZZ0SqHkxxQXN
DY8BD2vp5wA3ML3o8+hS6x35zl/zmD9iU/uJi3vYeaqUVumHfnhjhFAhbliPITaBiFW49exNgsNB
rfcfFi41aaroJybkkt8vNYSyhb0/fCiuOB6cwrk3rYDAwiLFf1uUHAPLb1Jh95x1Y9OwPe+yR4/w
JVN9AH44q1lONDFEbvIBSqXq6eKscerAnTTSoZWqfETOx7qdubgrwCxXD+ED007xvMFoVqsBbV0+
hZrexRTd9m8HAl9ToVE2lpIB5w4cVph/R5PauvaRidPvxt2/+SdLUxWsgn8RQ9/kwW+gFX4dlyNh
6gBEfttQD+Ak1mf09ICLVn8VA/EOE2uziRbzKP/8KIM973ihuru9dLgTkP5+pvbgA4jeTRX6Ik0M
argDtt7cK9BIp+oKo0HjZqyooxC1qmf79oFCt3zTtQGgCDafLMXN9s1Qh+GKhwCax5Cmerl2TZRm
4f+Pyjzgw1CyqfXxREOF0DXzN3UtmihO41ZnRVKNLfzyjdE4e8LCgSOA4SDpFsA7fGWmXf58kksV
b5vdPe+eGGoF0PVs39TgesdOWP2j7wB2MIphdT98D6xWujgJI3zfQOnv+CDQdpm2VgzWIeCnlybM
OMxWTKrYlJa+LhqAqF0n43vBC+LNwT/tZJ2aAelFlUizu0MsupHuCPS0HlhMG6GJuLcqzR0ZvdZI
DiVm3v44m3/7BmzuiBa9gr86UdR1bgKE7Yki/YSXBVWV6Wf5jOD6n4ZL5qbBIcasaDQAC/7oFH2J
bREq3nAOp3Et2JaFmGcgRpcuyLJf4GH2hEO/CrR4wKtRAjv17Abz3djCkxy+jQLSjO+7yG5tpoAZ
P/mvP8HeAqlJM88OH97q3Q9gDMxe7+Y7kH73Ew87d/WBBpqXqa3RNfLGtDxD1YEey0O7/lPlVx6u
mdKgfgUr+iB2wChkfdytpWh5gTXUr7BO2ud6GOvrPSWyhqOmg0a0UtPbjFDuWFNnN0uOy6qH2ta0
6sqcGibBw/urKpZTmrZQm3GoKTxuMAjY+/hDaHwk1oWU9+jzG0Yz67DxaqY/VVUeyi+Vo2doHQr0
b6dEvC6Bc8A+a538M5S6pYnFwPp0lLYHxFX1GaP3LXLttd7wyEJYTE/JO1EPgkBWMYO2ybb9v5MZ
oNb2UL6tACDXTWrOs7SX3ehsMnIYozvPSeUITg//jTkFpVkCk172vW6Zm1ymWmVHcwI8lhTpl8kB
xKNyDALUZ2k4RPMX6HQqsgfnhy2WfpG9tdE4LAHmYF1eAeInGnBsYIxNipkF4Kf2+Jx8PNRp6rhb
1uGq0VbASKsHMInL1G081CdlfKatBdpx4ljNzLHzC4UPK/EkMyoi+DldeVtM1qSUXXwWn3Gkh+pN
DSluUJ5mfsbx9KfQpcIJ49thWHd4OJKrb1OrFGZjhJbTPe593V1JVxs=
`pragma protect end_protected
