// Copyright (C) 1991-2014 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1.4
// ALTERA_TIMESTAMP:Thu Mar 13 15:23:41 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QFVv1yghCFIAtQ0nyQffwYU+hwfuYeWHQssOmGb3X+hSvV5sWMdmhS/jvCNl4zo8
a2EMTA30D7H1lmFsxSfh/UqRTHy6IL1Jd8i8JSCDYqXwKLbLuX28ybYhI8bZTj7a
NCEj4Cp0mOmzkSJuhxVr2JRWmBkWAoF+q48+1y90/nQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7488)
2pfcrdk5IfGJR4HiRBRzYsJS9RSs6gJFeBc4+JGt7yMD8c0FpcR+knRnl/6gltt4
P0ROcqJje79y/ih6c6iQRwmQm3ZWKlHtdq+Hm39oc3KCiO+TmOyGChyGvaWWbzOU
e6RCx9uea0XNdfikMyuBjoo3pl8eMPKgj8dLpP+8tyUUku7RK0lvHkt0mOPn7eny
FqcZ3YWCXgdXmKnFDwLDqq+hJytdSxmVZ2qTVLN1VOQIwDGGzcFXmRV/MrwJzQQa
R9/Gq9NNw3YmhuB84ARmzcaMNjPF+0D1NkfzGQ5a7d7FRhL4lvjRykbgvTUen+Dd
qIKIY6WZse9c6jZCQhDEUQHXUN+MrPKdmQkSVYaKEyXtTJuVJlHLJaXP+dUYTklt
H8+hVm2KFaXRhAj/ZUOwNZOyQlnIZNfL8jBTQWZy6UAMBl8ZMhf2JdSnnZdu7X8U
67tSL52X+JmaooswqmCN/t/ohhbm0lbkgKWtIsgUsNnc6IVRkUN/J/abb54zJ4/p
R0uBol2NB4aswNyobZcfi9IpyEc0cS6WXxGJDYibTUvnos5juPcoxyksG3n0rqTW
hdiAe1eKam4bGuF9T4dtEzX5NsLnWZpvNsAHO5zDVzm31zfD2phifyeV26oDcdyQ
Q5zj87AKgMxhD3FZoNmEfvTgT1h8KK/wX5MxUy6W20K7vZDGWn8+Ka6o6ceBCxmg
HY2Eact4wu0Zrnp8Wa722cx+XvzUyWX+rsGH0TUIWs7/MLXSPYC0YvSb40l2MmYc
O91JpBPfvp3FaUYtkHXE8zApa+BzobhnVQL5BAlV9RQuclzhquC3CIo2qTbRM8q3
PlSMWtJbXvLfBCUmI1juo88ytpmBWTwa0EXMwatABZFXaB7FMdPcV80MvHypG1JJ
E8yPZDXIdMj+dBTq9sdSy6pTK2TTGVj8rwBPVvPuOU8pSnXwW/7it/wksS1RBGNF
16+bw2H7JN8yDL10EyP9v2sV4jFjy98pq/syMzeu57Sh8zX/4BN8NPH9PojLG7tf
LIFuam77cz/o8ViTInBhmc1xbY2LR1tLwhoznEDwi0JTc6ES4bYYl2q/XlXL4L9M
gQDNyqT1zpSB8WyLqQFfjR8+MQtl4hXWzIjDs9tdPkDU2tPV6Gr46yL8m/veL/p+
CgAWwBLZz29WN5+vUZWCVXxsPmRq7H4hYXkjUlgU5gVOSpOIqvDibvZJqRfE2nYl
+sRIxu9H95PlYkYKHTAF93OzMBeN7bzU7VkrSxNF5MJTNWJxv0mq8ehYdYCG2L2X
p4F0xjJEPdLaNlxml+sWhYg/SSIZ3Swo8Lom/ILF23sg3uphFudBRT0Oy0yEsH0P
0A7f81HQWsR49y2KDtaPfy1PXNa9WEETgtkgtGqWi/HgfV1Y1d/BVcrsoD22L7Gy
ZOoUm/GJyl2phvDtyis1ivtGADzCnlWd2HwAIqhXaqyB4WVGbM1qxiCPOv/oMkIz
JmRnkoey6WaGUWdkvkkFkXLcjwhn33lP9G7jnWWyexXvfXiiyfOYA1y5LNDc8QFy
6x4sjipwIK1aEy7fekrwyWMk6NMYwPXA2/8zOxEZ3wxXTbWUL1kxTGR36qSHAm66
IiUgyjLEcpGYAXhOitRf+2q8ek7b8Avc0snHYosAtyVgTSJpUjI2Lsw8InV6Zu84
MmfGjvBKIH4dqb26zUHtvHz/O9uCGO+4HylUF2U0rv0l4KoXP0TTUO+nfnzzT+6/
7qLBxjOt9JwlinxDa2mbOtUgPVMlWn0pw3fvvwuaf8i2YtgXoEEjaeKWUUFjps1+
tjNb05OIuQyLnQMjtL6QB2N8jbtDBWK3LGqoM3oKZuzYDc8Chu4o27EoY+86slya
SZW+WNM2DRVEho2n/cVKHh/qfoCHs7aQSJaAqioCpWHiws5Wo98Dqkz5h7bm/O1a
RwsU/uCqsHeeuiTLESjfI5y/82CS9lk+SYh1YYiM3e6htnpUon5OWsKz7U3ijZgr
JmaRjtqP+umw3FmME7GDq1RACw6jeeLin2fsXBiND8JH/Fge1rTT5ceOGbftjvCv
PKpW0fVENxBkmrTjFjOf5xf+69vQMms30vJ23GCSmUr+rGzv/47jLPJwMoRi2VNB
HeP39C6rwPrDB6nUp6TN5SZv+HOUeGqCoc74dXemsXNzdr4Ep4/AU9nPzjOLmp3n
CGWN2CSontuMWsk5lRJ4C0sykcO5gKvRDTve6I/318ZG71KpoKiAQhri5oKh8ImY
aIFZ4q0yZXUeWs7s23mHrBnwPNHx4seCJxbGSWf36V7dz6RkQtvws6WgoiLOl2Vv
cnLf0s66jiCl7iyNY2g1VH89OByrM/Z1ICdCOLiAAY+Y+58uwEg9W35HcT3ubG8b
yrhgNn7052IxfoeBcOk6iz4u9Z5TLyeIqVWKeBSgSZQMmsy6ZB1ag6x7yRM+uRSA
nLjZWt6C9t97Mpv+do6sumeKLi12+NjemuZMJ9OcaBgttAejlK1UnKYELQcAjEA9
BUOUwXwiCO2l2PIb6rXdiL6280atqQ76Hv37ckFbi0YJojjWEipHUQR0aeQNMbpF
R8945ax91kFZdxJlSWt43q8ygt6CVIawR3Pp+m3hkNvh/SnJfPbgzPiBiutuZf/O
AfB95wwmFHmrMQHGZWsyuGPS2fVLW6ZW88bMDleU+8BX8jqaUPc2t0axUUvvx349
jxS+2PslVVDH1+HPzjpktGIPH/X+WrTvXoYUGIIKADIErKN8yQdLNLsp1laxI+Ck
3hQa1kIDHk2fIdaiZn3SpmUJaj3mF3QI81/VpxtbPPHheEio3sBKxYUC7mDAmHWe
KGTGEX28KDDY9Asd25jG2fW9gFj+kjvDb40PjrHIOUIJfUWFzMZ0rO/IPvJzSHBa
PDgEosXNI7sTarWQVujsxh+ap0c63yY495t55oXMNGkAEciIsV+Lh2P71D/0Dl1B
aLifXA0/tTbHlwCQ3Ry1gss6A/WpYNBObTmCUXl/O6ErghOMh+kmn4F10CIlMyjN
iAj3U9A56lnFlCgaImXw6Hkf4Xcm4RA/KS458hoozq8GPBESErK8ROblljVWD8p2
LDrgI8zhOZBD9WGeyD2Uv49ux0i3Couv9sm+JN6jQWgZZ1vPf/nRyW92pUnbXS32
8G398rtVxfP42DeHkFJPsA22ECVyU5gXw4CRGnurttW9TTtFMInCuz0yrG1K8TOM
epq9TaY7nZUUXTvyrVT21b1sXXdakdNKl9Do5mFVPpCikgSVyB97MDddT2IWSM79
A6vIXmk596c0GqsrJkiXwXz4D9wH+6I+KvQSDwYGiAOlqZ5KeE+qP7w/4KMp27jf
beVHdsn1X59VpNCofnS+GcthcqlDWPrNG9E4FICC49nbt+z6kz+6NlA4mdXy+4pG
xAUYv7msmO32z9PDCxXXk7pJhnJ8dXNWilk383oe4bM8JP+6QFlA/BOAS0UP2oQQ
KSMN7ZlCAOhWmtxZkp3pAtWP2AfGky5J9wPsbKwYUFI0SyRpibS4mgwcA0zmIxaG
PTFdKW8V9PT3oddv+jWZA2HFt4gtJXxJdo/fNLwGmvqHMfHZ1D87ds/aNYFaqBQr
cIbCzT6AMRyRfSgfcD8af3Saj1VC8SnZgPJovdQTOIhO7jB7lA23nABRN+LnQ+VS
8XgIZ9EJ3laKxvj1dUfzPuRSnp4CzAmT+sc1J/0xTlIBMsn0Xg2hDCzqWPE7DHu6
X86tR1OvFTrkZ2Z5G5+mNm/8FyZDNrRfoNCLR4OpysLAL+L9dqJirmFANB5ruxr5
uf07yRfssw7R1UD7sdcXixL6WryxEP06Yb9MhAfBp1S5r8NZ5bz50ixYc63gqIBo
IQIkYA5ODDJhc0DIXNungPV3elpTFARMlDDzjXCtFfLkD9cKKfN7pcWMSqHJossh
GxcdVk/DRcFN1vCZp4dWjymnUvy3V1r6dn3FTn7/5y5VStqqxfD5VXSzbZfAwhqF
shakCd3YoMEjTfbdNRYFw05V3xQu94z4BfF79/GNOmd1huQM5qPOUGJESwBMhvcp
imikpcp2FhOWh8bQOShzdtnkh10bl1UemitA9EynKdrDxVV9dLaON6hGdyB7tDkA
al8DazK2oCX5+WvoMBbMfVXCav4teOtGqPesvzrKZElTITyqqIPD53+dTBxAjA3B
WXhFnEOCBVmFTVUx4UE0csLCctGUyCSGcoV+ui0qzjXSkXkPLFwHV+dd0l9MOn1U
elm8DU/CqeEWOm5QOFqVfh4FnfFd5BplY5tDGXdtV74APY7cdqJ9815LU8NQS9mi
f8IkgDPWCR82QoUTZYmf4s1dKAW2w4s6fKV+peyHS3qKUewHwwbnAkyfnGdEq7Wt
nAw0g/Tdc04iUJHu+ndlbO2VfKXYZIeYLjOrtD1sknOP92HNT3qCW1LPNZc1aqBE
kxCE2z87dn7OLH90yu7fp2+a1I9smtEn2uFwj5LTw2X7AuqMsGV8SJVbWIZ34yQS
8hur/fIat7lhy7Ru+sCenzOEReJhqQr0zBjaq1PZY7+rYMOvcSwQlHsh4a1p6HqB
J8bjxpLa2VdTZdyeyavjFPr9pX7JVlIcwsUapVowwG8xrmooLG+JGZcbdtBcrVXC
YwoD8vo6c5SY5ODX5kb7ynIulsf7i+lHcc/G+VJPUqJSQSW86WYetpAYftUUSNrV
eEcJ2G6dHaPr8VSRFghrNPrOb0Ww0/LHRaEPXS6juwLIDHmhD8lNAH5AhSppe2Rp
SqO+xICd/KL2aofsd/CEMYfP1tN6j3tG/fs5IpS3QoiAeBMQEXvi7qpIrHwlDyDY
S0hVU1VLgqJ+lxI5BEMv/4rhGXL75EZ0pfWxojOpeAoMzjp3DW8XsKe1i6PfAqc4
x4nwdqoHyej/lP4hWkaRO8ro4V+K8EK7eExOlYC5WBI3EGSG8ITKzJfBfkCPyHT4
SA/G00KZl3gAIvaiXHyFQYJvYA2uR0WyyFbc+hg8X4e62UENkjYHcq5Oe7Unevv0
hrNeUUdXx1StgahvoiqA2/rQDAZvdLmeEBDV0kZdFgP7oCZg87DfLaGmUqmpXFxm
kIaXRqoc0wrsU28IPFMAf6o8M+PIn5wG/ZCzOHK8yOofhl0/hR/rDhLoIb2U3bxU
5n6E+U3VSgvxpwp9rG3vaYGwyyq9Sc95pAi9n4ngCigUrrxqDbab0rWGpuslnp+w
/mNX7DS037J9Dme49CydPtp7OQ0op1q2TaSC3oyGDOapH3t4PvH9EUin508aXfu4
ccffCmTk5/SvQx6u/mAgZmXZujF+a7K6dKhSGfauz/8YISGt/UtUipVpilJOfl8X
7siyqnST9zfpWF+makysjBJN9OS9PLUrWa+nTaOgn6zoBklZYZVJyySGS84aRfgX
D0CxxD05W5ISzX4OoPWsTXT8gd9X+KbPxf6eni4dN7qEa1kglRDbPoac9E2z8Qnl
MjwOdtXeFdgcK83RWnmfNymNJW0weBkFTMwmAFqTmW+N90E+9LdCVHjOTgI/EqNk
XRUtX2DvR74QuyCSWhWzAhq+/inGRhq23fW9OuaWkSMWcxeZXoCGwJdn9q7hVEY7
jZ0nOpeA8VYu0crXkSItCbx5xwn8VS9KxUJail50AYW+6mi6oayUX9naTIAk1WWR
vXbH5sI8lhKHxA0/kZu4LwDgxYC3rEY3Jk88r62GN9evpGmP3EQJbHSFoz0uu4a2
ARWqo7eDg0mqFXoJn0aDMKT93yv+K4AVpd5N/hW3iGkXvBL7mA4qB/+fr9eW+2qQ
LBJuv02N1uKQKsV5yulpLRWYb6t+MvSkoBYU8p2qCZcRzDTdlHyWte9ZRegKwI/0
uoyGXHHnud2W+lCCJQnxwv1PRS8WmXYKUFcmvSM3OSjxWc88LXYKd60X8Bt/+u2+
RXoK2g+5zWIePzpXGqQWyy0VRr/F7EmPS201qkjLSfKPCBOtOtTKeV/u14utl/wo
8gr2S5aWFL5pLb+P+DfYjUeo84sT6CGH2IHUTLfJlTlwmd/A0yUYO2GMzba0eq2l
sc/uzh+W3hvlOAqENDfNnwd7JzhMkgKoflpOifsj2LgHl0R2WSAPlj2KkxPJd0YA
exUmDkD0EZNo/aXkuF+IMDwBdBqT4gpljZ/J1BubsZFR39+v0steRhmf1cmgY+pp
5KdAz8dBHsN002PvFqBvknuBIPqx+vYbgiLK5IV+EEj/RBRC4xE7P3FcoVqN7/iW
uLM71Da+qpRTnA2iEF0yXkiQfyoLLXb5lUY5quAmnSacJsl2CFYpHY4q85D9GAP8
JFTbd+qT+oSCDw0DNVkGsb1lpaLi9hj6PjjBso6u6gkrj1u1JUMnMpVaod13tuAm
R3YrzYvsygDEtWp3ztV+Pm1qHswXmHnACqjWcS4MVj6/jGF+OgtCbJvBatEGGCJk
vVB/CqCg5+rK+YrDvuj7miiI4doJUVzPSPf4K8npQv+WgcDLhLoP+Udjifv6Yp9d
Z0xffTP8DZnYhkyN114v6cQSE7d+5QJ1M/5kLtFx+dg9fW5WjVhRmCUD4IerO1yP
N62LYNbS7vmQuvtx2WLtL/hyoH9qrq8xMomdT3eLB4KPdBiAopKoueZYXSxQEqLF
roEGPtBnA5WQqEmJjrbCZK2idrBfZ9QUi5ubFmq/zIyVxt2J8mW6m5dkd6pmEC6b
U7jet/5qzVQb/76fHE4E+dg66+xlFNWnhlbOfB5GXB0p7GTeKyhB55Ob42Oh2RIm
3xXh55ipZ9VjntZZgf8Z9skRoF4uarAi3xvbQMJo7Bq9EHXBqwx57XajmS6iUmFV
8P4LFqX7qOsVwRMHVpgb1BAmvsgTdx0IjoSS2/ZQ0v5T0+ofViaCi4zu0Y1jz/zU
5/d79r/VFUXoS0dbiNw29UHYH5hFRunJ+JF4RMPCq0rxbHW4RgBfScflHp2YYVkB
+DYhls2XJcSs0wGKxsymDI2ndAeG0GVkXulv023wR1UtjjBYqUHxMCPxwi9i20zn
Cb2su8LSHgq4tDljX7z2XuuAc8L+6SRAepaBAB9JMN3tvDMgA74vj2CyfdMub3A8
YTFpptaQfQk0vZfOILcO2jgXZsTAH6fXtyuz+S1Jf3o33CY8Wbll0VSGuVv9WXbq
4gTdYG3JzdjhK1D4memwZHCNLJjaM4naUPNaNXUhB8xOqvj9B2hOIM82/usM8r2h
kYswevLLHiuA+Cw7eR6hXj1igZrW6E/vgGShZDYqbQnJagJ+nA/NU/rG0tR5VHjD
40A8Y7xr7P6lf0X2f2JNCMWf4XcntgxVZQkGSAhoE9Ne/MWxylkELZcPjaNtG6dv
GD4ubdwO7CMpzuuQePu+fD5SiGhjyvLOSOyKTAHH0lvC5mV9i0ssgTiH7/wCAxqL
+xjTZRM3WU5NNugvAf4pyFPq3+8uNAHveq3pDeISZXJ6Yl5vxboDarnpoSjuFyFy
OIzINdlSpg5xJeX6CDYzIYpGBSA8Hs1POWS1Pi+6ylLwE3qD+0oeEgUTTUKcXt9D
6FKPpeYA440W9+jzJLXKxSeipw3BZd1Z2acF1sI+sNS/FZ7iKk5TKNFixHPJA/WW
iW0qOlxJhJONA4Zx8QQ1HEj/GBTAL0yq5pC1+nEbemE2tiMXyQTBHypEXe/Udv4J
pCIuEbceOJHKYYwQzBr8IZxMd6Fl8RcFWKDDtkkG0xU+C7wE2P7xFERsg2TS8UlI
0X63267DPUQVtj5gOBh+/MkP3NR5saP5CKwIYUS/jF0aOd/KEisokxqZMcGaDAuP
dGhwZJVV1JUwlZlPKH+gmHBsBMObMv2bXZXjhBtHj7ZgqLMrMogKQ6o+habjA2Cg
Co1MPm5mpx7I+ZYRFB6TR/0bfzuFXbSgus6P6agRhXcObxHGu6IEWcm3hT6Xlhdl
lJw/qglrGsymOwr3/+ZVTr3jtangXKLh7Djs+nm2yUiQQU0nr6saMCIPPUu81hla
QZ4+h0nsC5Ugm0ihuzc8eo4Nog+mX9SCEPLoBKJjV7tjlgAqKQVGbGvNQq+sod4b
PvAr3Q0MwJ/FDca0bZclfXPSvoev2HzT/K5hEOWpSoRmKgpzKfkJMxcp4sJewuz2
RgIIv/ewO/tFZGpO01Wzc71iyCa661b40eHOUDNMdg9jMOh02X6gvhS499p1UDdu
CLhEjAN91/0RSDp18KNYK3tXYEx8yOIqSdstTHLdc1CRkVgPoUp7xj5xQCj475ta
Qcm6k+I3eTaozDHTDb1mKDVbA8qe9ZWQNlZNjT5T6NMIAJknNkYZz8UySsEONGKD
v5G6oww+5msJnxtf4EzS6wN9cLlLypGEd1wD4srQcWNl+qx8ZGZ93cM5D+tce14m
F+RqPmP8YitTj+cFsYqEMfVLatBZSinu+j01O39Z7PNlCKk+CGHTthcyN8JLvzhV
vKEPzlRuqn3cfsPr02uEbO+POn1PDAJsgorLKeYaN/PlYS3SLVO2KmwEzOES5DVn
OwAbx0vFTwHddubdArAdAxsDyMDN9ZGQiNvb+GxrzG2cyt2mxuLisUG/MpQRVZ06
QTl9ZgUBWqzsJn/cfQZXcTvxLIPF+uwTTi/FTMwRMKm9hHbP9V31F5y/MlK40aef
e9lgrds7UfAVnLGufI2gInNI/dq/DvWB2OgilyzdEou6LLpkMCYKmGNcpM/2Ptrj
NHAuFOdtXDlqT9hnTa0k/Ktfc90ONy9LuClAfxYaR0DQrP6O8UbwJeWbGJIEx/2D
PWu2FCgbKNoZFKNuCEm3hkNfgQPIrK7aE0oU10/FDbm4qvaXTqw1+iZSUGsYlbDP
JynF2BQiWYAY6V1x+rzWnOVhX4EzwsfWC+wNKCMzrv3KXY8nt/Y/4/ZGKdOksIaS
cFex3QLoFHAnjzfk5JN6uaU9EdrSxjeS0HdFUXYHbSKFyZRbLVFn5VKNpo8yjQSE
L/arfsFTECVigrXSSkC25Pj7lFXIL9FQbgvGa32oA9/+f2oDTaPkDZtn4KVkgaxd
PQRZuiEcbSdg0khyQjW4aqYbO77tVU3I/LTCh5GO1YIYMWVbsYq4EVpLq4XnYtNJ
j2GVCxdF5z1tCeyCbhVgjJ+cOcJHkeZCfTfapc7sXOQYJ16u5Q83IPzONcqIjcLR
SKxniBSazd3uX/8J++qIDk7ThPZrcAeeDcSgyPLtGmS0529/aT4JZfvMcUdpPkbu
lNDctL7AwNQJ2QpNbau8H1IncJahLkzAMAcenmzC+OKm+pIxdvOTBDpqoc1rG5et
w42RrqbMb2+iwg4IFiztcaSZAbiTNh6hQ2fLwMkajVIZtrttrmsGiByOEPCvzspH
qD3xmPV4yidAZ3glqOsTR8VFTa+PoZ/ZVF/YPOHYmnTzZrsLAOqKEXZH+3rBc4n6
ZPYkNOLotXXsYfBu4r4wFaQ5xN2Xs5QbPbq+SkvY4JTBNZnQXwBswW08aobRsBGx
CIfzc1L2jZP59gCOXbaamnNIbximpKbDwNJiYOyaeW6eFCx3lQUjpH5pIpHvTcwZ
a6Kx7mjR8ckEXgI1BybUv9PwDG1OQYcJV31jemaHcFQZgqNgRJeFXWTtXKWyFrFH
UfmkE4QbRXcwZOiY3qPcTGScHhoHnjGWiVdWdvsTEbJJrEk1czAJx6b1CPWkALzn
GEbmvd+mDXRBgaOt5Rjw17JDbY+OdgkWVTbIG5SojnIiOLL88Ivd4JAPZGUcB3/i
RlTeAWRLjLm7MoaVhfoYBT1/HTA84m8ggrgMAkKB0L3iE6F+rwFbY6sB5wOcSBC4
FCLyGOyHkIgHa+XZO9g3utwhNvkS3TWPYBG8lIm/oMCpfZ/yCojUtEIm5hWi6UdA
dlM+7AXs8bnHFIURg5U2hrFuJnfeSRhcR13cRE1jMRMyrvYHluo+3GmyB9gGDKcG
RnHcQFbXGqtxb+lv1qWIuPzfIKMScgzIZluaX5BYPHQvadKPoTy86/o8+VwClkrw
kkr8hPVxGQutbHUyQicpUxL/1rlZ5nUjxvPFULuDX9KQIUlhUSe7MdDhC1YeZjL1
`pragma protect end_protected
