// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Z0T4HDLLrsI33sqikk0nWdca6s5exi3YYceY+hlcqxVM6uZWJu28zk9Y4OXfEVvjHxCGu/nCIJdG
aR/+8VC507PiTvAVdP67OWOwp+dpBDsa98ron3MFkVcvTknK4VtRdE3P93/3hZyvs/OSTA3AU1wW
BLJ6kigq5RmSZPAWigT5PWC85olEq2IVzCrkLaa+47uQiKNFoIYvlqMW8S8OqCqeHiA7bGRkNCQv
Q1enxES9GCPPzXOU1HoiuFPIPSAPC13SDfXMH1wRE6R+cKKkzlwGyCtRjdgjfQ5RSU2dHCGxZvNH
42sIMXFb4vUKxMuOmyttaqNS/ymlVOkAT2Xp/w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
kuDz6XCnetixAfZPnRWpM+Kv4bK3gVx0Wl+vV8XnGNIjM84xQ+l0gC8iPLZSK6C93FHEm4zLszUC
QzMMXsGtQOQERRXma7RbcIWWLvSRYDEjr2SFB3Exz5zXjlqmDsaqo4Nj0b7NYOo3Z0jYZlLknWPd
/MXdxcU9bBDo//CExmrPuxMNvmOSZnKW+7e2UHasAePdeAF4NGNC+YPWNSaMWW1q9XdkQw6Qt0Zm
/ME07lPtYxwjwL6VpRINDXJv8XT8eOa3g1zY0kb+ZMIERQ/5zZg325N8pnAbswHynWm9U1/0/hUu
2j3tyLyPwp7hEHgGj0TUfo9tBKhae5+orMXk8/U9pEUO/VA9J7d1kTtmV6oF61+E5eyz8LTv9gpd
5GVve/WgezPMRCms3YpkJPIQgTUB6a4RbkONNDXgcQCFb9P8p5JDSsEuzCmgZAQk9Ej6kbfAPwCU
piS9G9QQ74Hgu9fzhW7247eMrZ3LwOR31p8u3ecyYpJ/adO6yutBt/Mk81pfqIHJfS7jtVHa3/DO
ETy2vnvCpVKCIXh5mcMQYJjK7z9+gM6mt6BuOvB/egqcE73M5AHNZXeQKJzyozP288Z1AIBRaPJX
m3MwVLtxmxCMGK/Y2EFtDm8uRcuRCImoPPi6wfdQOrpefNVpvgJyyu9hrfBc05BlbFglFL1d9rXo
By8jfcJ8FMy0hSG7DBQckiSo/+LIapAp6FLh1A2sVpTwVgPPgeww473WepyILY8CsQ21jq4ca9kX
CDEZ0sz7Pe8/nZpr7maC+GrIgW+UyOdKXhym0wF5OlktTNmZWd6orNcL5XnovoArZSXrS6BKUAyV
w7KROMah4H0eiCUL65zT3YziXTGLh/eZU3bwQaB6JAKyXFoOwEJCyqWiqzFi1dRNPK+LLOS00w7f
c2ovvalCrPOdelwgQWPU1exUoc+jiwOHIWtXEwQkQBPojbpCqEecaWAvLi2nR/eJeNhm3lL3gvP8
ecmo/jat1N4K9SVyIHARD8KZUcqwH1i/GyrUQ6VfL2/fHSfJfrG0bAy5EiS9IOqOpolPPqzwQjGE
rtRuhIA0pV1XRUk+Y87zSgcOf6RlElnPbNV4EhBq2IhWhQyvJixTqlJeo2rVAF1b13whUylyYrAb
GCQL49mQAM5vsb4rXx0bAwJBxHBrWjg8M8p1Y//vNTELPoB5ZVrWU7A76Ay3t41hJCODlqXtneyX
ok/+5WHJfP1tMoPzLbbzST8AzJQlhi5FPVc8+9dEj0WRXmanPLGtxZx5sho+f5TGERSLMGTI+Kjg
pJ8XdWpdtH+Sz87wZvp3C4EJ4psbYOPVXmpsOrvjeQt7EdctgXXC5bZ/fZ0YuFdA03iz8FtdD4/L
7T6xr+O0US2EiJ6XUl0WUuVjL8nKtnUFk1lhl28hSP5gIj5H8n/B3MuoH/3Dn2fE8h9AKpDBI4H1
628tvmgcT078v4GdD/2NFGs3zPKmVwfYhkqo6vi8ZesbSUefxI2Nj/y0+gKdD73Thr8OW/apQZH9
C/XrWtJsiP0CggPabmga47v7o0duqLOOePh6f6PRTfZ399TqqggT67VN1+Sxh6ATimldZNyz0NiS
jtU/bo6/bpAoiE89cwMbEC0i7fGbuYS9eZ9GNKQL9WOnWc154qMqrOqtGi+9V5fFfBh1GDfBaHGW
mincJrb8MMv+AJlZNCVaflbokRr7zUfNf9VXq701VoaCPihibzRwyhllNJf8hEKzHJOYYGQ4twk/
Tj9kC9ATWNG8f0SuYkL0D0vicBxBX8Xh5XIycWzhHXS831RLm+ZwnjDQvslSOeyWbdSRZ/SVrlci
oAQe6bKhqerPPOLNBTCi1CJ+rzbkRidKFwAtdosuxBIpBz9LkQ0cJwALdgUhsIMavVb3pRv8eEc9
FOyirk++jGTgUPAV1rRoUbelT+E10/ldIyk9iH64R2XcXHou3aCLTw19dQvu/kpoO4XJk1i/skLC
QHYFG7J5SEXfotAZpwZkdmpFh+mZmITbtp1/QqA2pDmvfTZCUfTxGh3JbLaTCQZC/gnn+VysXw8S
qqx6HHUfPRk9UNPArYHZHJz6xY4v3IYsn2n5syt+8J1waDDKUKtQajVDtI6oeRruCibhom03pc9t
P0U8hpsxl5Kp8qVeqarW+dJyLuxFRUB7uvFs3oRYJmdgK/3jNCNPiQrOu2/aRgVlfjClf17Siz/Y
zu+WM6VNI5Ure92KjxXs5oASvO6zrOkxt9L1+LwexIentdkc6H6W9l/2HZ0/14XICMFM6DS507O4
oZJ/UYOPOAR+Namw37GLmwG/yGHmPBeWuv1bG4OFOUX2frh6qTWqcl9ZSeKRv3SEUyexIwbiaSyx
3UlzSzhG1Kq8dTn9m600to2kpQIRQyujBy8i8Af2ZxMI4+VPiYRaxPlYEfRttx4IUUi8tSV/d+lY
jfaCr2VryhMRgVzQ5a/NXUnzCvvqS+mQvHS0b0iXQBhJYJNjlBqr5RFbrS0SemkzgoESnMhqHXyF
5saKo/vcL1Du1LkmrB7GBbheIxr5weSgnVHQgXSOKmMRuN4+YGN+FxdTcp3tz/5ubNGHddYlhzLs
KYh11ROGa4s6Ckg/7qaWOk5obMe4dNeNEHC8SzWjtX+Tz4LQtYwpvn53cCD3RIP7zf9Cooqgt+09
e7XJjJxERvCcwqdh4bZAhCUZ8glBImyNyBFIefYLOPM68YDUvlB+Bb2fbPB9IPDxFBMzqbD0euvR
0yOYpe0XrXMFx84kzv7WrJOwB8DfI35XJoeunjZOnXGedbKTcTCzmU80O7mTBMxoDJz9aRVeMrzO
wuf1FeYirfb44L7WcVgGsoTqGsCws3uV0Ua1PNySFl1MQ6Z4/UlOU4Aki5iLZcXr4xdRshcQUtK2
G8It0/nLvzG6KaIkdwhakMKULwvo6n2heMbQ80IvbNU9RuWV3182fMvvC+ldr/+h8aiHGOqeSb/+
+jVk9I9h9EhMOWrwwQ+ZT3jN1mu1kwQB3PzYNCJqCDhCLG9gbXSCWPnDUhsltCaQ1jQrAJbF2pPo
bNooFgmKPX5BGFhktF1E5ofANKCGq7vgZ184mC7vyXENr8w9wVAHCho5L15rsfFoSuTE59bdjDYI
ZeJt2OZ9Xk7Df7nWqgO8VHDDbQ3kE+Jf7sAhCF2fPGpP5kWAPk8dfN4LeClQeqLcYogvVwaVBkr0
aKRNTEd06GhcODSSnbjKHAv8sb/9GfjcchOkdW0UCjYCixEPEb6yOSRkC24+hMPO97W7+90OFuYY
9IZ+8fmNXtMLT7nH0/0c4WL6efm6+WBLXKnbxJzAedXILfA4ovdegtUqb7ZE61ooes9Wx+YbBoet
o7cuhu4Lye/Z5FwxHYMSX9gMJzwqFCIuCUl8VRZaREgJEkcNI/SpSPWiJCvBIo/66GIihkY98zYH
jFt2ev9C3lQ1ECdqKppzqPzgHzoG+dUKzRKY592I0lzdYtA7goHPBlioOKUyr/uIE1H2BrisC1/e
5FpSAMMFMO6RSqvf2adU1iLGsY1cTV1hCbLlMKE5ADJzKF6/yAhjCzvAB5efFyw2dmoRlWVF0KFH
64GJkJTBsYRq5MhvP4Mp2J6+YfzAyuzFQCtdc1PhG8RuAF/duAuF8qKADt7lGIGDSBdSa1OEpxpX
KFfZwMCFPM+2huK6n4gNIVygalvnp6IuLCHz93ddfYqUjQCWWRZvS4WUq65QtjdlP4WDp+wH4yET
73s8lYt8DqsH8i3TYlIDVJYTnYEYwrxcqFsZaqdnbl+wjBtV7YJ1mRVYlZQR5O1LKVoX5t2wH1D0
Ug+J7SOMZLUBPhsMS7SKc3MtMGb7aRAThDH0dZOgbrxAWtUsyScKZzBX3Om0W3TwQiisdvJUWCgX
hU2q+Nc7rMtCWw/wefXJaBSoYyNL9btQyo+M2br+9z8PGVDs523VrKY9c6b+I6HH6UqYc92N+hpM
wUaf2Aj2KA1NIEtzUDirRrt2pb2RuwgEoqr2mPXzvZZidyhuSxEwQw7Yl6afIOaejqZLLQMrfBnV
P4P+l7nCixTs3o+K75jO6Ggn1D4sMB/cbP04msYzbTEZKT6WcoaIr4T7z31V0+EvQF/u17hToXRM
CU0D8syvA5mrZFilbl7UKeaIU71deHRqNd4UgEFMCa+OKysydvM5rdeciTXN/7I2SL8x7FzSI/g6
dHDFcmp22xNk6mQhk5p49zwzJT9/ZqFswJWbO18EsJ8jZS5GSEDriuv6lKoMZxpdXmU4GH126/cO
K+9VbHEslHkArUYXebx6U/7208limqSNaouW/6zdECZuwowm4GXYlOE46CB+tVIYdmatOI+6zuNX
0djcjP/IrDVrWO5WxufEDS3yzZtvZly6N5aeTvIx/sdUfTnwf9DMAEvPzVsI5f3VawLFy6cbF6NE
OuyOjkgQC56ZmLHOXK2MIBKEyieCypQRu36EXuVWVVbc5jQ1zouAvDog+sQUpgtFS7ed+UJt8wHR
xsbcQjnpTsaLF8tQ9bTHrAFvld2cXUkreIjIawh+jKVsZfFxqQtqetQgTpvkZcXDd3X5kpgDNSGW
kQKKf+wJps/JnaYuNYW2E0ccV9Tv5ecEXFFpnuy206p9wxk3RxXfXh7RTtstNP2z5Tzt/8YpFsv0
R6lCLn6TVFSgTKqb9HwQ7qTrd/8giFFIvZ9NyM42VFbyiMShzIUvBnPhxr7mksGTciFeGDiKvuNJ
bSb1Ai9mKiL7SdWD3Ge2AoHPfmbcU3NRS/5kPVQiN3vobYOE7+MOn8tloRGcfdRCSxLotGTQPnap
YRNbonVkHSmY8OMwuFRcSDzXJVJqM7Tpe821paVUmqaRkea+WwFujloEh9UKaKlAqrQWOgH+ulpL
swl36PXRKpBG1Rv8Myk2RiCKs5RbXwnj/UoO+4nopYApUO0K4IwmO8Jd+uXF7Cna8MSrWT8+CSaY
3wGyacECTOnmgCw1TQG/oC7h8X/wAfnIVuX5yVXl5JM4ezPo4ylm8/lOo4yNHsVASssa2oKUkncV
+rlc0y+jKPlsm6OXbzwF3kgp6ookptbrZEK+yrgh6kr3MDMe/EUugT0cupJXAT5svpi0uGiMolFY
XeZ32qGs6K5YWVsGZlxbOGgj9fo1D0XKO3Pr5CZ5Y4d678mWFTGlX2k5q9hw5Xmm0FbQBGxRkavp
Lqa8rTP2/oEjOs9MEHozDhEOwnNABPiWaEu5b6ZN55xN1HMW/PrQW1frLz/YFplBhO5Yo70Swx0z
AJGm5FUsY8Mnxj1Lbtdb08fSaffPmyNGfKLnnCLZc2Lw/tmEfXE5hbcqKyw9/Mkd5D6gjrF90wwD
qchaMmTlFPaPZnev7GUFIQWkeQH/6E/cSkM4ZZj0OeEA8nyImaDIDVbTl33tf2j3eX9rtRbcAnnG
cNHVFBCZnGgkXk60L4Uf9MXJdLw0CIYhSXFOddiHM9CLczajS214TyRj2wT2YAFtaDIJ+XMg020m
GLW3zqhhcZbkwC0IyJor3dRedjRDkp0l5bI6gcp3yde1NNoEfbRWJq2Ra6Rl7X5N/xzT4V9QV8cK
/jQNAeN/eKA+N4bihANBjz4eSg4gwxoxQSG4tsENJyfR9zxLj60YbPPA+Y7U6g0ZMssrQsuebFK6
yUELUlyl7tIJnOd4+YhPbSqutvUxXR+pF3SRFO//gKnk2j+vhYWPVCrt3k6Gc7jI9LxPa3dKBtRk
uNI0RDKssiSV81QTB7B1fx+wVdZnBgqIh2ae6XnDl57z5JDr7fG12iHDJEZUyKCfANUFixNQ9qpt
l+t6TN/zcog+5m3UrgcOHebWPE89SSiE2C0BGug8JtP5CEHtJLc8yvebYYy6QZoFrgJJB2/79etB
xq8uSSAM7DjaTqCef7809NBoPcT15lOG6gO6SiyyQczFIvHHXiQY5q0E92anzUm9DFPJhki82Tex
yJVm2Zsa0YyYpvo+i20VljgPD7AG4saCXyU021GfOMFe5bdT/gvOIppFBoG4DiiMCUK7J1yhdwnN
zekfYumoTZizPRTb6AAipdDl8doqXCZFX7YQ1YLDY1OXwD4qL7nKGzkoo064+RWMahv5xn6TFLEi
h52RM008k6n6BS7XVwCMweXstNmyLUBmYb15BNKIXrUY7EaNuQd6N6ZEka3ulzhTGE9XqJkACnZl
w1r7wDWySaF5jP4BlUMJBCzyMvwDEWAxR6Mfcfqnxp/b5DsAKWT6gA2uR/H9ZGFPEMeCZAKCMi9T
+tvpZIFc82Qe0yFenoleAOBYxN3HkZ4gAT5aYlU9j0Z+NYZ8hJgWTUww18dK5IG2KIKfx8RHjT6i
wAwuSj63bZ4AD/58SvHhWwNZePnn2G3pZuhLBEMfAVPAvX21nSp+87KDam2PKbbclIsFD/IZjacI
gGvCA9McK3L9XnXXSc3axEyMmFFt4UYBJRwmNv+uNBb2NUAsLYoOTYxA2NpbY5n10jBk1Fg1OGjX
qpPTXjVfq0swkTqhcqPPu/38TvI0N3nJ+/obOJ7P/ae9Orm8Nsb4gRWjLzP/Tk5YAGTOgUpLTnkE
jPRWo6VO19SeYnu3rnGDEOEqe85OoNWt3boiyKvrfQ9aOMWM/EhAFEbXcGLeliX+wPwvoIzQqRKJ
8Cdn4vn+w8jwGYooBXoqv2/j+UQiEATn/ZDQqRRslrpnCPqfeSJCRmh0jdmq+3bsjpOeUc4ps0S2
wK9cb49GZIvcaJiRUkeL+9Bs+bYtwsGVQ//45IRQOOcKtIXZfdSMPAlqFq7Rp3/u/THKzJLD8LRr
7XWKymfaZwOhpW+11UmHpJZ6QLLdmR5hto2VDvWDT1SZu29tVoZwraccvlilNvOu71w/hpz4kQ2R
Yqb6nga/ilidfbW88R5xERGK9bfZnFuTHhiajgAEihfpBq7iCzAA2fygpPprdoiM73qgA4P/ibtq
V6ihq8ejiJdTPEPd/fqVBEvuiedaO7mr7+jC1yZwTjbizwJnZPG2VfiF7X3uQ5xyi3uF6LiBg5E7
WtAiYRnMhG60OJylZvNvcYlHrGYWtypJsId7riQO/hW7IPnlZ24vVOGNqWDHuYmi2wcIX654A4ZT
QbnbR1AAAJU1mmTdP0mWjfi5/5y4MpfeIiocN1qA/9Csuq7JaVvzNSavH8JySM59u9JE8/otFlFK
6Fjl07DKQvEG7uH7CMlxBJiLSpIHAvAPwVP1xuiqnkyQxV+q67R65buxoC4PbUWmkHiGr7Zn0alB
iG6b6RI9FIVNqnvkBGjLHC312BuBrRXLHOiUk1oUreU0IQBEXp7RweQKY/w3TiTrVTWSCZOSQuta
g1MhsEs2aE+qG713AnlXULfFisdYN4qSOSYrQeR5FIGq3i70tZ1Px0IbjqBNzzukoszQwjRDBKFI
x2BujgIoIFWczbqmqq+IpKpXKMg8w+R+pF/xDLkUyCnsNelsai9dv6nGXZe6H5XgPjT1SwEekil8
Azt3P4kuc5ml1KIWMwl0Rm8HvqltLGOPV1zCFPIOTMIeOZfVegGkfdYAWy6kcBT/RsT+nWhYKjd3
GJhOr9L/3RGfU35wQQIYJMG5I7lGdUDHkhWhESfmAtCiuEhNnF645Owrotd4gN5qmzI908oCt9HS
V+qNJPPb2SdV/JfQTo1ofFRDi1aynv6xwwvXfBqFO2BKhIE3lS3CckOuMwxw7XCFiICoq4aG6bTj
WCy25s17DXkfR7xWEmCunf191LqystNJvTkj4sJpg89C+ONFSJT9VYqBuCg5VPEgqg9BaX5g6M1V
5XuKcVYUYNcJAp1nC5lR39aXRS2nPnDn6YIB9VEd1ojWslDbOs326Qm/gwLnJvLlUPqxA9D+hkcF
9kd9MIgda0am//ykehNcsorpWwDRSw272qEo2KuHvEeUpve55zwYSEeZshEioaYdy2ZHWnotmvVQ
7l8TZBDzoyTSQz3McxirX9cco3RaJz/q8Fmm0dI4bWZ+lclK7gP+dhidjFpNW1UGzV80lWc7m+t/
lbNPdlRLQRFEZ5PrtNYYqsp6CiLIFnhU6VoALoYHXp5olnXNaB0gyrNYtOftaZViV8lCcuQ53R63
b0/xC69QIVpom+Kq7dorvetX26Osj56cJuPRfFUbYINdNwz8dam1dQmJiguL/Ch4ZQP2dg5sZG4j
LYk02o9bUHkUevGlvXSI+FpCkMUb8cRMK6fyefPCNrWhHQnE2YDJYdwCGJImmt0u/KDs3dr/zKxx
Amzh8ZEkN9XOkdpuedaTYf3dkFczLoWfgjpYYx3MnHIGmg5mVW8iRTkjHA8vgfoLlx34v4arPAM8
wpb8tt4B4VZyXxAMFfOIG5jms3vCcWdPO/3OjDuy+SJu8TNTcgv+R/I8hnlySaIDzfwP1dRUW/BG
ssHvmb4+5bYGRS8yNfj/BI2i4ZGsiQIq+F3/lrNxlHbeb5VmuWwWm6loenEyWkHlJJcmu67xebEu
X0yeevm49WlJDh9HHmBhyOlwWzlA8i5MkAe3JCGXGqUNm+XIBKbyJO84FhJFEweq4fN914CMFlMb
6W33jZeglhBE3ivAlxIv/j7JYQp/FZycEuQnU/b/Yf6GijN1AF7zecsQI8UPkmawGjUlwd1it7zT
fM9DqLvzBPE9tx4if/HSyiMXXx2YvzOT170BHX0thxO4QmSgUmv7OApcBPEhKza6V6kJRgn3NyH+
egPzp5fafqRfEPCjrzFyhZfEY8ujz+YxhlgBGfZTnYAv5NiDADh8l41G0JR628CQZEoHtEK33KZt
kLJh2GrPVWmKz1yqdhbiVPP4LkVSLuTKnU/E3SqYXzrcGkHKjrn/EqYp863lsbHaXrR4KhgxNO+z
Jb5rB5ZCQdX8SgcgkuZ1f4pu4K/mPx7BuuK/Xi0/o0bsxf9QOZXVtCr9/7BDfikNxSD/SuC9a6tW
YwtPTF01u5BQFGzp2UZVl2LsUKVnT7v50pW6NspHpw1Wd4Dzevno9Ox9Tl8MOHK9LhmOJhjDOAWh
UN8C20DYN/IfaFzLXcmjl8IPr1YD6D4m2bCF8NKE0vOLs6uU462bvtiKViSh4mAIy10RNuK8nQP7
uFEzaqc+FNFP+Yz1YioC70aRvh/pCId4PZlNaYWxsiypGO77e3NGyrbzVKk9L1fykyd1vOC0V31n
bMuRTqutgq8C/CeOyRF+dP7X/v9uj943Sw20jvXoZcjwBpNdDBu1aMRi26tskXmM9+5svM1owozN
dnLsc+6rQo4kE7ktLZ+E201ywFQO7t6S9VO4ywPyLUFoEpJC5/1/YQ7WOPBUKVGxT9Tml+YQQEvo
/tgOaaHMw4AknHFyt7rOBwdTH9KL84fhsmf69RowuTG86RmNk0eAIgMHCou0+guutO5emEwTCkoI
B0SJvtUvvm7A6PS+E4GvnWyb7xc2ZnyY2DNRnAVP1ZyyT2758HME6vgkh83eU51jGsRk0bHahGwk
tfiR2a96Pwi2JnGIqiLloKa0jmsnUqwCY3szbLwSp2j/D/ko3WxuDWs+zoCGBm+krdfLB312qzod
LYbzTxQXcD89ZXZUTeaJNahky7tF1EgcCUSY+4trnRt6fGtNKzPuT20l+GA1756o+0r/6cP4mNqk
aBd4VG8pw0Hy5ubLYkm7Vp/Ki9ForKReiWTpfxHJMm63GlhN6rc4UMlUX2JX3RAtnZNAxBDgvfdB
85wwe/g9dA3ZBGI02W72/qFBqgIBazZhKH7pE+xn8ukUZ0VhIs3V+NztKmu0Mew6M5s5X0Knzoqx
1EwZttOyWQFms6zB6+9KiSmLugwmbPlcTTt6SQb9Kgd3aJuETUbirdfQs1cTFBS4LP/lTuqnbZCK
BxmGNUaBxZhzD5ias6ObvriCqtsILzKdVFe64aBPScZXvQUHhbGeN2I4SBf+HsIaOjgsz0S3ErWH
KmjtfNq4hRMfaTU7VAzOmHHEVzG6sKIClSKsg95T9pT5p/d7gfk+wAhwYimaXDW1cryBq308DKdp
tt/PsRLaiot9rmRcsO0avHx3fJzNKaBDtdsJovkmnU4QFfEfpvQNg87YbnI89isfJyo6GBB3GRG0
glEH6YjeHIAkYmjcANKZzD9GSsoVK6b1ULTi+gVrPNIAIZV3TCKE0X8GzEYNDdmFVd2dunCt/lQb
hE+FnX6XMpR6AtiVBmtTqpZN/MYAskRfc6mQQxpPMY54YAz5Bi2fgeuD8rzP+moSXx0hbrkAJq1I
uMO5SIqbmuxNLiEtYwlKFht4KjjfMV5vHpHWhu0NQ15NsElBHKuKRl5jh5yFPvtaZFVqe1S7biqe
VEjFe08goNW0gd5L98PMmRqJlu73B1y43nXaRgHEkOmvpw28B93eEKYSgluNboa3Qc55jv35ZPa+
aTulA06OIxY3fhYjdalpRq+fpAqEGtSAS+w7UBOx9C2RK6nfesmiIYgVP/imnG2Hyd9pSiQlOaw8
tZWHTIUSFndUz0xz6Rgdco4xZ1uNL2Pnq6m9yLDkdms8TmUw5FcXakWWZARYnxMqmmi3d0hontEi
KUDTxKnirhGOk+6MjEqwqEcZf4sfB8Kq+bYDt7tRULtm4rko8+JIHR/azxcH2iL5s+gJOblW7HoY
koK0yCfvKFlowW9qleIO0SIE00O+UXBXCO+K8ahLIvseXjvMpPtSHjJK6rKb6s3wc/2w8ymMkT4v
2atOjfSJGjujgIiGM4BqOxgQle/qEFzp5hP7i5h7dVklk7KSaRqpbZVMze3LJsnpVDKJhIRZiNhD
skJUc1yQ/+fWtVp3sHHTNb40buH4CLDzfNnbxwi0IZcOJ0yVfJu9mauq77c68dUqJeyw1m5Co6Tf
GHHS7oefxF2e9ZlCEtGjEX+CB4yLBD1ZS8pvpjroD3fPrhHwoAHSQshUDWSo/cWGR0liJ7yFbKh9
AbN+hvUPPsIGjjTCOSVJuWXfPKn7i7kpR3yOor44FWoA5CweVTenb9WBAPyQ9NzHi19ORufv7imC
D9Q75lKWC7wkFbrJk+4WHpKrg0XKrhlcIH5Wj0k4S2mu7HtJDcC5j4gX5Lp6lud6A11EOfVWKZjY
ZYSR0FalXz2Vq6UwkkncOMtmmHVvTs8cmsM3CYHJlMh8AJMvoE8pT9ZlLhEziTCpBUVWj2vGv0EQ
JBW5ILvXokTycE9stK2kPymdBjEHZssQBEdY/T7J9UekRA/EW/fmguKS+OKi4wzKu+V4sbV1jg7f
t92/atfZ2aOUIrg+PziqdPN/mRa1Xphp6zkC/DPUt54d4WN0Gb66Y2OOUciPgyJrnH/Uj7piEFKV
Tuco5mJJiEgAyOGZ0BSsQ205t/gjvb1e3zwCsoEKx4IPjY2GAwdg87en5w2Oza4wHSNJEfIzd0pJ
cCusc9Jn5NnPPODfA/q1neW0Iw9s6vRO8DnQhQnAbCzln/Tm07GOddigyToytBhWE9n02PZx8qMB
RCmAiYcPugeJnv0v+FACu1kKP+PaAsWrlKNk5sMqztCkExgw5wBqU1ukMMCqlHu38zvI17+11p4k
Da3M77VHGP2NWaODADVdk7kX3Up+OjT3IzE2+Kq+OSLj/tjEgD/pw+NbJQGU2VtEmKPCmEovz2Yq
TX/rW7DqedlrW7iYnryucxH/nIkKR8pfWjJ9rjN1+m9xHsOwkiX+N5Q/KGgzXU5OsCEsHHGsYPoI
1c8OgXV4powAFNgJH9qFGEjR5I90nfA96+gCtwOX5Lk5BC8ustpoVhgkqWBfjdX2fHkr/FVN8w0e
pOnwhrhlX9v6BxhBBUPV2jrXouHjyrm8/RAFp+XzNSmMQDZm0AUqs8LCQkqiLIByzD0ApRXuzIJ0
t1IWUp5rLjPpMpeolhYAutJW1r1+vWy8aUyH+5eUKvQw7E1OOomdkLO3SRVgsl7gAqNz5qBdQFfq
+hCURLO5igspJIjjJKcD7vhi3rYYbhDUgKNsScHGNbzMARjijj9KPfXwrvCADTUVI+5HMH+USIIq
w0XD/H9DJzzh2QLbSe//TbMBCydDrErBS+KoEUHd8Vf3Ivy6ksBvyHY7f7d84yXp3BUOO07naRm2
Pe2WfkazSqezI8bGUYN0JSb87h4bRVA2UwzDYXBWHeQCgPjJHxqG4z6pDNQWLnwCDYlBLA4GDypO
LaaYcJDioXkGf/fdMAyXJVkUqN8iSSCJYA0TjsdBDuiC4P1vLJs46dJ7dmA+TjAKemmBj/hfG1SF
NfPcNNinQai2/3Vbsu0M6lICqbC8DqtsdDABhQ4GsTGCzE0zL961lZ9rpj8cOnbcDlRN0j04ED9j
h/Aiby+Bj7vJ60EgsW961+cVJCJZAv2eWx8GGv9RO1iaFlArX7MBRFQxNN4xHjUSfv9BkDyEK9gd
2ulMInpkVy6hojLUxbDr9Uw6XM01V/ZwYwsaZrAymXBXt+044bpU2WeKJCKAjRtFgBUa+gmVaEFs
Suj+C+L2Q4qDvcMZPYaqVhYnmRm+6AIZKdTE8RjyUEepxVfOVl6Vx3FIj7aRolXVCRs50bFJjT0v
UwJApQBg1qstm4d9abnrrNUGZpLJn0xBqbuoG02Jvdszpg5BUPoau8KWjGzE9tN+cwx9bR/RxL85
HTlw9JgRuYAg8kHoQazBn8PFklTxoH1dv2aGkQpB6dQ62fyczCsHpXJcVCnI1qI2psQE
`pragma protect end_protected
