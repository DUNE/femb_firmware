// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:51:51 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UT31HhJNo6DMB5GVcqGlpBd+cSXsIh0Gxhxza/VI2phUjFhgkmBc0Sq8yefTzayl
mZEZGBLHb0vwLfnNz54w68qhIaeht9OWZxsaC+gEU7vpl7k/uzCRWMvieh+cl8CU
fcM+h6tlcIRsczLXbXHO+o7gOoxtVaRdjzPz0sxfYqQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9536)
zqACeJ06wUMRJXzq+TSnEIw1pUPpkcQ+AKsbw5a5mSS9xBgTMIfRjf5LV7OtCDAv
Sww/jxi9I++AohDpI8j+63ow060H7QTXH0Y/Z0t4PUQWj2FEO1IxySmSQuv+EWys
THZVEtww0hURKH2ihTbhlTDCOtgK6Ujz30Dzh6NSlo4dcfGz4xXfC+BtFZ7RsdC6
aW7jjlgxt+G2TWKsDROlBmBBGd6HaNub8mjb7H7ObhqVA7ZFU+eZbEUrVAH8dCgB
lGGkrfPl5sMhJpmMQDHt+T4NSoLaNRxEw6q6bxUZrr7qdLOmFwN1Stm0phU8bOOk
cScxUOAOv9VZ7fdCCf0lp7sJR4ZX9ArhScP0R+sDKMXUjQ14COfYv+dql9ISSKen
2PsYZH/u4ITXQqO2Nt2cjP8AGRGkg0ttayrwDe+zJ9QgSFu6Ig54j0fI7ZlykJfJ
mkLDJsCunQhUTiVOJPCS8B2cBK/MgGWM9V4aiVSuReOduQYHvSQ5zjSKBgtKnQ4d
jvBygrgqWiUwr3JFbBuNlmR2hVGoZWlYm+zmFKU54bLww0M2HuglYDiWCVjRZ5u4
N6KpBT5EE7ZkRiM0QnPHRj4mbIJ1iY2IOoGdwamuKl17TdrDyyl+Ca39hIowiV3p
K73CQe8I7H8NMogqvTD1jqfgvX3aU91m365SojYa/qrQOPBCb4dxBo/81+KqFT9q
HPLG2TGAex1+NNtV9qiR3ukFLDeK8Ru7lNbNHFbmdV8rh1QjqVpW9/wiVVi4w322
1HYIX1dLyW7tZk/0Hr/XPaWOmQI/Tj6cMjvCzjUR8jiJALohWZki1iDC1Cc/Vanb
+xvT46f7kx07c1EbClL74U+vCXHFIxM19GDo5kTOOt5VAQdQoYjIAjZNxKJXLqHy
yTwSaYxiW6gI63W93D7OjXjyO4vPKq7cUgt047sHZcUwyIl5tRyRiMIWCiracD7U
YVO6u762vVIXto/sVo6k82ngF2lsnh5PFfKyt+g/x3xStgjFmNhPlTD+HmiCtpi9
an2NvWniA9IysTzB5CKDR8pyaEUAskisuNK6x59IlhNpxCU/ccwgQhP1Ah3+wmoh
beJ6KVx3DyYCJXG1dsawqxTo98n7RnW8YMxQwOfdFrU9W/V5tzSmtgpYxliZXyIy
YUcjSxrpzMwEkiaw1zzvArLGrjabroYlq68Ob323eWrcjUqj+W0O3GFcja7GiEtW
DDHeE008rKSe7IfIcpUMO+4dbC99ZKCYHoX66vWJFCuof5oPqPcHvfK7ayEMXjC3
KwCMhoosR+s/r/MdN/x4o6cDCJ+V2jI6fX61l4owOg508jTO679sfTqW3OG2QZwH
x/N85A90TjKj5L6CMyQ2SmV/WVkKoDDF/Ey+hdxEHW2grHssobOsInB/F/35/aVe
zxQsyHC1yCqphVvUxco7as5zEjpLOahV0bnFWJftmPzKOON5FdpEDsL99PcPmzOq
n0WIz1EwyzA1k23snkf9u1eJezSVY1JuExGDM5px7jdfGYfu8jh7VRzoaA/BsFyr
1v1lke+8eou0oD3cBf+3ejbrWNdw7vbzrkd8vS9axsiLMFczbfHsUL3AY2Wyg0ij
WyZ8K+KVNAMSF7zulZ1SwSKCOm0oqRzkdSO7O26fTc0JYLTEMEsXp/TH3q2r0WDX
Bqczl7mKgReJY+7LA/qGiG+bGv0WK62i3pJScS3bSOc/bJN0a0LKHHOD+3gh87zt
fe+mISbgNH5rNGablDskdkfYsvgihUarBHrJji1eZyIRAvmZeay60I4GwG36qwvU
9eWuW0v2VricNKq+gfPHhs3x0SGA99Pr5nJGx0Ofuo6Fqt+rOQSMl/r/oTqUi4rM
/4OyghQ1dOmy/4klhsFVWybhfPkm1Q8BrJoyV1NhzHRjZA/O7vmQ49DckWgYszZz
+VjyJKeo4XX/ERTqCm1nLjEkPJXFMMoIJQpQeBstkSbH6y8mp8IwbIZ5dA5Q95LX
Ke/QBJKdKasrGyze4fmOqEjo1rAyM1c5gwEkMWTv91z4bWisNU3oeBBwusPN3jmF
9CiA+cQ9eL4tdkdXc2N0reDO4g4yF3Cz0d4OiF2CiZoqbexmLNVZ72b9Ka6IWNP0
cGyTenrU9FVUQhPtEIeQMbu3wz3/+EnSmKQ0lkN1itijt4vBnT9uxju37R+QrC/z
0POXuh6/t7gHTDXHOB9LDBlWMxAefAeIKPKVk/7rDPx/6oMgUXMvPdiPwLA2SOyD
hHLg1MvlBRAm2AUf6KhlWvehQU1x6TTRreoPdMDO15afu4fObrSsfBtuR1J30pf3
r6T9ht2oi/UbjDJbRQpOyRlB40LGA6bH5rPO59VZbrDiR0+Bb/Xv9jpjW6ackgtk
f3K3gt/MtPP55zaT228+hH0KzXdNHfjP1ioCcIUmJQkWY45KCYN0B4PFkmi9sWGs
2icnwZvNR77DPrpE37oj4iyO5NOH4dryKypW6gLeTGPyRm32VnxGrOWd5EZffcIH
UbZPAlhrAx3dIXPwn4eHW8A8s/LqQkhbbK1GZ65BJ9vw+Ga8LF59fieSbT/zUi/k
RjtCxLzbofD4fQ+emiEOElrS+4VZ2PznZrSZvUCIphp7gvFyoC1hN6se5aBET/5+
KKqvsEtEjp8Wyc2q3zn4zkGauT5LjAKu1MWKFsMRmKmV/c9XzEgnnsTaSITe9No+
9SWTgJvcdz6Itr78G08lP2tjmDp2XJrk8ekZ4sy2RwO9yI6yMYJlfc6LCSB4nDJI
UrKZz0drKPqpqTsh1H+SG163nYUO3ijrdfjwYrsmwACHzBUeRi/abkYPQ295Hlrc
KdSgX1azmqOmoGvAIUNew4WwbFmTlhYVb86UmpGfLbsoiEBxuSFMoW8BeIFDPWYR
cIBTVHxka70fLBVDwy9MI7LLfEtoGlA0NkcwerK2C488oU6Ohc/XMNgGpWFENyox
ggEqUFA5XQEhCkxX+A97/fThg6IOWvalJbSnuUUy2HaKP9I5SOgn6pfg7vssYNtO
UUKNe329LJPcUjzqAY+xdlLFEcvoQ4LxeB5sifN6zTTNuHpk0SuF4449JnU8uj6W
Z2XirfWeSNz/dRBL5+pdKaOZMc3d7Gr0lieupjgx9fJBwxnbRYSPNOKDMMHURhQC
kR+WZaQXi0DS+yfxOHDEBDjYYI4buot4JT7bodrr9SMmPbd+zHPIgn6JmgLN7exi
ViAb5HzzLkPpMCe+VyarNdxIkEo70N8NG+SF+/lnJH16tMWikpD6azGUHJgH7FYG
PNrkQCknFO3NHIkLZ/9OegD1z031JAJcfx9RG3yBU5iqySO0VkdWwk6BaPuIoxBX
2J+pWKtGO1cZS8piXJ7tU7xPRB2h0qNQjLF7cMf7Mu6NpoV3EkowGurFyEyEgfec
y85Sy0jh7i40ND+ZG88bEdj5en6Ps4hKMDoaKf29uJR06Nst4mHRUwBfmR2SS983
h/wWUm5WUWpiY70ZCt1dFAbVah5a8tfXJqCZyLiEcZR9te6n1hnc3isrLAlHarr9
Z7QLYRQ06c89LaUhM+fSwLHjycbhHOunGPnWgNBEseoCUs1VzF3muIUQ+ai3DZUz
JVSLBzg3sIhHzYsvncuAYwq9Y04ykHrk5ktSmWNb92OE5mO/G1MJHxc1ZcveyU2C
S0wgcmSGxLMQK53bPLYly5RglDzD6obAqCZaKACPTwFTkfwZYZVDYRMKoIq8T5bn
LhLtr1WavQjZjUmFoovosqEbL3I6Ill4fvDwqFlolcYfXNQ6fXV3PdHtDLHPTdXs
BV6iCjiqK8hc7uH9LWK3W83FR5wgNpBwjNk6upfrES2cNDUnCzMC83y8pD88Uwyl
jM8ip/2c2gR/HcZtGOHmAJeRnkD6VHlyoKCjrDCrtvycAjNEMauFwXOBTctleoLP
gh1hf0bYa1JIJI8TQJR0Yrb0SEaTr6FRjsMm/mfyPhFFL9sLSis+wGv1B4Edx4E2
Dve0FSX9PAzk6akmDi3sIlcJ5zpjzVATRlhG4mRL4mX+Pbm23HicJnODH2FOvXqN
+dHUQtTNfCgU+zFBp97doS4CNOaXFq3ziuIIHx771iJeL/ICa9q6gWbS6vg2sMcv
GPfmX1sUA02RTSVZ5Iyy1MSzblbfq4bsenNg+x3eESMLEIFHKWgHUUW8pmb1QILh
YtV8P8zww1kLoxTEiq7Nuenl+aSyNfCI6fBjCBkGH/fgCj/cTelJSTptGiXaDbpF
H2krNA0beyIMq0NOuI0pKGCT4q5G8pjZNpc5h3jGr6HjBROC9QHwPrpdqEKQIhIW
j04RV6u5V4d2bCCbqs9cDQpYAyDjI2fap/PbJI6SVGHnBSeds/6PWgi138JkTuhz
43bWS79wxAQpyKh+pSRH6AS9z5bFST/TGjVelHjaQcYJSk/t3Gfm5FXQkWd31E+3
686PW12U/OUVkstBTwyb0QTvKZEenCq+b6VrlnBw1c6lv+IKQPAkeX3DkLPE7qck
oRUIFTvSJf0qPT/dZ627TvpKPwGdGMbLTt8ocVYTRbWYK3YwcZ2D/Y7SedlZrwbQ
VMsWnnYestXKy8fmdVG4TSEkTECJpTBq+5/XKOqtbeOCUkcJr2wYD5WDoTUQbNKh
mQyVJULrTE1HbbdZluiHMYQI85DUwKzF/cT1kfrBx5l1J/TTb38PsyazC8VaVkOn
eCtsC0nouTu76PkfAO7OtsWHgph/t3vo7GIcNIhgiIFIkQhtvpXuAUjtdFnj4iA+
y8obYH0wWofP0bynWO03S7pAEdu+CMLncHc7nDB5gthq4AN3f5bAlQ0tEAVBDbLz
oRMNtkSwZS9LU1iDTGDwGI2ehToPanKb4EihPecLJ3N1IhFSw06Df9lWJKni0i4j
6UlT4FEkbWGFY9w3w9e+7sY0yBF5vCBUWFCCfE5+aLU7i10aXiyhrvHyl0uJcNFj
KdIEfONF4y6rs0nuPz2VEmV2y2l4fQsUntYG05qYFTwze9DtKGP9/OzrUYY8Vt1p
GuF2vQm4iHlYtDIXTy7p6PV3D/RGdKIvf9t1GPTwcW0ylKEezjyRnBKchvZf1j/P
PqaWcLamjEQRONwRRiTxSSEFT4zKW59VU0d7ifKQ1rlUY9Fy4zR6aKDBe+6yzHAF
foukZnwzP4HkJN7KrHK4sHwk9A9hZZuoCN5oUjAqvGmFLx6+6cHWGMDWh2ooS/i5
QK8NuQWSLaxNEcqQ3UTK4pknxBVw+uqJqPiilQpndepNiXCaMf7lvN7sXFkXwjQW
3b1UMI7lZxPlWaD6mC11WGwg2fjHs1f2XNz625haXjlXFojD/vryFdEwato5sZV8
stoUr5EQQ159yGNkq9u47p6DhVKD4wKl9Q+/XZ1KrWyb89DIKwPQGY83DNVcvb14
ALtSnUAQKCchlIpPTp+7wuZqKmgJhYHDrnr5adE4qlUf4dGnRVnui4ELT/WXPji/
dRHJMBc04JLb1UuziGXhSSMvsB3IPG4WesHmrpmvbBs7zShFpM/XBenBff5591v0
/qMCpnmhuxbzHbvSXWb+/UAMESCbOXVv23FD/QMEqFhHAaQbYjDn1MR3ElwsZeTW
Z7oR6cxiDt3AWPCEBWtyhyet3AbuWZffGTNW2heY+paTxuTXO5GDoXMIkLyD2VS6
eAMsPKMqz38T8C3QEEENewNVPtXgphU4v8+haigvIxo33b6eqEoXRVa+s1kqR1yq
Pw9/YQrd9phQ+nQwG/fzNBmQCPh7LnO9/5Wf17GIHw25Fd2P/ThOz00fF58NjFnK
4BbkgjrLAgXVRk4D87jD3SaAls7LobpP+wSrJ0GuLHqFshY4ZrgesUSZ2WwvstMZ
NnWw1WoBa+uOEvGuvM780y34fQ8nZrkAB4r42nfnsI59mB0P2JAA/husjbUww/Pe
1bsstY0mPqV+5ZlJ46tQqtPXU8upCp3juIJJ5hSDonjmmyeS17uinvP9CGngGyII
Vbh4LtLYbcamrz2VVqzVqzYJzl3fbPhwzZXwuGQ03C1KFcegkTUtBF6LIGYglJy7
7pH6h87P1LjrkuXlaIIZSu3A82fbwrB9yyLUt60WXFiJX/Q/27571pB0C9NHP6UV
ICNVVOQviLcfE48bFoWmcs5CWy2mvb32ZfPqA0QGnjbvxgs2bmcrTu9rzsxO9xRp
29l9qyD6pCS4iKZ++lQXul0IxmqBakHFMAqKcVGR/f28WftHZzmhV2sVxII6C2Fu
67bVr8kWxFSvKywTpT4x/FznHtsi88Srdp+UZUsCYWVmny16+TBvtbu9nr8Cn+E4
nnOH3/CRKbXJUNnk9weVNeWKFhrcPZI6UTCLVSRYGpSG3b8Ny7LJVXUVFbEgz7+9
xnpIjsspcY61odcCRQVRBU2gL4DO3+bB4mGGYHVgW1VdccsfxNVtHgHkb+bkalLi
HsFZyxtLT92QaAt4hMQyvYTZq09iJaXmnfUg/SmMpfFZWjh3QNJb/3RiahxInHiC
T86G5M1eLP743s3NpkgAT8VIlDSo+kA92JYyb8z7szs6h2qHWP+C163O54g93auY
O+wGN9o6jM+Er25TBRSiHVxQMqLA/N0pJg2KBMiOINNA8nCOXBd1xYi+Pm/mRzFD
xK0Uv8pe92UupXwrw9Xrqcpk7M05YWrFGuJC88fmPHyLhG++pvc3izI1UvXOkn/N
mO0m82Inrc5dAf/8/ZlwlUAQxsqDSrQQ+IoOAb56ZiYAn0/iQDBJHVsYx6/EON57
HGbciaLG3FgcEI7loeQrx354d/AhKozQ73fRXn4QHmEs4ml4FPiYvV28LqS5DuzZ
oOMxzutRdUJD1KLHBDuqK4f/HjmipzA/eWYyxoTSytnBgxCY3LOOpbZC7MT/s7IJ
HqQDjl4LLbQtgJ0i/xQ0gf4md5MLFeg4rxzcV6E51qMVcyCaIPS3CIWb5RD/Svih
y3MrDMF46+5diVJBl7m+oKBZUL186GP2YMFqkfDGuy91P1tZNgU2NkLBVK9gy8rv
AvUpvzQKbUrqmEpDH6QYhbQSQzmurVHJvty45vLQW2Y5erDzQcBYmz4614ABBUOx
LZhLly8HxP7SWGmHraj6ToyDhTVayilxPhOYtQ5W1CUM6Hucl0D1xqryvB9fachE
ZV5AlJq4lcwCYiDfMB49nGFEq6DWHUxx4wihc5vo0kBC1aNMBpvhrXLAi/FpUUDu
wpe3h7cPcJ2csrjYSVrUm7NwpTgBNEWVLq0D7HahAVw8cd+waqTJZFsNj/cOgAuk
ZTRcbIvDVbqr6WrdKo3jULSDSzR7FUR7mMmo8D0bzdql0wchSv9UeMTDiwsHLdEa
XOFKaRO83sJwE2xcRKi1DzBiiI/pC5KPPatVFXTctPLUxJGeHBoA4wfQ8kttdWOv
gibPJLngucvCr9FctYPnZSf0BZEvuU0KluTDa4WFpaJWWmcpdKukg98x8EJw4Edk
uLfPkyKYo3D24PbRTf9LLjDUVvhIyXE2YZTYuKGVoSDNRAllnBshfVy0kQ+UOoxA
GgI0HdoEBQE0fTqtJQmH1YqfqyNOaFruC6LVBXkHw1sGPmHsP8BdgBdAEgxZZ9gX
liInQADVAXanC/JenHjEEFixwUFJM+sDholn98aYGbA5rmFXA6GnmKRKw6EW9D0c
beer8G9dCTM4KEVi46mbJskEWO9CzPlT/bYuWPwaQiQV66A8PP0L9KID5STLKmGt
Ec+IuoCj+hukjfqz+F9WOMEb/4zUqFi5AvfjIQwubDHcjN7GHi1J7mKXNuXdeRmk
TNc8Ev99144vTD9I5epgHPKED8eb6ezhEuyjQJQeWsLa3XvhfCi8zCxHLELUfOgR
yJp/7hDXCeo2lRGp5rV/Yl1//aW9J+6/E8pmLP72kP2SFzoFslElywVeh0GNuzDz
h51Pnh2ABGWMUYp7s8ObEp+cJ+e8DkW6IJ0dYuv2L0oyQPMHxrUX9sphTrI75T3W
Lqcp2d1ZTTquHHMzs5EPdKuNdEVIfs+JoJezhpjVxLNqk9RDpYRj2JJSAsSbBaeY
u0SrX2yYnKNBIabhCohCyC9fyg6FtL0MemaY7Jtc6AeiGN6hfn14i9OuUg7Y7iMb
NMxIkl1tDq3E7fEtZgbtDzivre4bwxVt8sCQWo2Ny64nq5QURLzsJoOepWnVritZ
f/rS9njKP4dw94/imHTvKoEYGj6a1xKkowH6SdFkkz9lfglkcKKHTP2bVmUs2vbh
E9cYJYEsQviqlUcx6JtlICifwtYlprSKZZeus57wSAFrsRHHaAcWqZUKdXxDhAvM
blhdiZ0lGP8GNWhJd5zVMQ701fmQoTn0QE8cDswYzRQ5wiU6KFGKUsVZcYZnLbFY
Oa8t1pCWmPcGv03oJDLYCE5KakMueKxub4DAjJgOiJFp7xEfxqUbdM5pYPkA8av0
4JTJ2yV3KzlM3tcnYjzJBb9c0jSDvMTR84VwjzUkacUw4MuwyPXB/hU0uGdR/NqC
oJcywBWua7mVlSvYvIS44YLQM5+Z1k7LEJfrZe51g659U4HS5YBa53TA/sYogBcp
s7xAO0R/3UwvJDUHriGOoSW4s+lqD8Nes35lU8GHx/FVGkEcEHHfuS4rGbJo/Kn7
1U9TtkYpVeCWhcyj2TouYBx8a1MMpq7sQKB/r7M4P0NQ9isSDSZm5FJWaCv7VIk9
8JLxPkC0ysXwqtzqbev04PW1DnhmisytcvovuUCKeFbweNZjUk9BGfI5KAMtt3VT
M77StPMm4TeniGcniCNnarFlNJm+Ov4xzWu3tB+TD8huqs4S7vntIapiu3k6bunt
qp1I6qrf1C5C2xoxjMOpl7cfvZUIMsbmQN5VGkyEpANvdVLkxtZzx791kWomIesT
+uIuDSOHKMT5hrwvxgTgwsXi1Hh8JC3q3cUwyoVpQtlgLuKFwhvgthdXmLi699Q2
XhFl1aA5sgAIy8TQzslhkkMoPZP6lHNfZEJL+TJZmM1IPvwaECwb/E7kzSASPlFk
PhGl8eGxArJNxPXGDxDZNEJOmYmUeAJerTuvJsWYjcpFkeLvuAeVMTEB24pRyERC
mFw6ll1dw9BgfywN7w4l7S/r9s2LTm+75z12m/jK8G7jsmgb8lkRJGYmCo6bxnIr
b6fueDB5pniErWwRVejZGVCeFmImlnvrZsmaagpUIr3Wr5TdoJJYZwYenCfhjTJa
RF8D2gH8GnE/ADx54Cl7+Jye2Kia6nHH+sprJLWNVaGXB/1fatYj/m9uHy1ReMFq
3Exq2BEZSlTfwRdd92q9el4K3DZhLxbznOYYWfiMBQmCMZd+z/8+3JZPvBUrW+u+
8QQAdw1pS3P/sJF5P4D0U+a6LazDSLBFeVvn7GdG4hGVdcsZutU/0XBC1sOhoD6U
E1puQj1DOZDcZeFzJQTgSbaGU5DLlI/lorcgVkD4jOoFi+3nBlCM6eGl8vlQ8/Bi
DA6/9djZVjjeHmN+UqxnvszJlVSroBm4Mm5DOH6lcLFuaiWDhGtgVOQYct/WHEYK
z8SO1x6qJU1w5ma4web4+5JtrJrTmQ9ptomRAfkLC9YUGq1bNcS/hnTNZP4vgXbk
UAq3QfsGJLOFFgsDrEcjhHMEABr7WkK+S7ZJHek8OqW56x7jASzMiaIk/O5r9orm
EeG7LrgQvxdm9hotcKRvxwhoSoJTiXzEYKeE8eVw19bAvkK9CTXb7XT2Q990BkxG
BlhM27l9TK38pyzrCF6BGxiusI03BzJmPO2KlONy5HjXyu2kRKublJTpXs8abJvk
LPt7SC+tXoUJAkWFHPZMuumVOgk6y6aRdtCatvT7PrlTrpt7R/j7VVq2J5+KyGRe
ATS24dTayl/P2Q1HqMySm92O3BAdcAIL241U+SsNZ1cSB3AY/DPP55KdbdfAjVve
48XDFcutXqqfMqm4FqN+SYhWfrKAtQmteFl6hFXTaS8/TBuuLKKXUPmZ0yOrYS7Y
/zjorb6uzEYsoPXhL4A2+pzVJlUmLsPIru41wDC5egD8xQ7dSvoQNRkYIkqXVZco
QB2LOxo2Zq3LKATUwLnrM1lTKVIPyNWo+BCtLNLNeFFxGG0puXcN/eoy02Y98AHs
8HT67TxyVEoI8ybA8AqXZOeLPa6zUcVJkfgzBxOnb9VAuJKRMJapsG0//8Jb6dK3
MKFI0yD03ANC7vA/ooCq+RrwAiCqUKbuHb4LjfpNZ7DY5sZnegX4OLW+txOC4RKc
TfmKudRy8NSKGciYQO8oGjhGrdMMzvySNBRApcNbh8DNX+FaWDdgRIfnkwfdFTT+
96OTUsXP/RAGPBtM+3cZHjQXgCj+vvQvEFT7+Xzm9yU0bOD/L5uAtO2MASxVVLmo
BkHNoed4kqJTaoo+Mqy+DEQ99Ly4tFAFgB8gCGcGvfB4SwqV2/JcnR7v4akdOwTu
0tCJAOOIWGnnIgyxKZN7ByV4YtLSe68t86iv1sI5WnQ99NsjlIzvjLXgrxJoecsq
aHyAE7L9qfT53QAhJYSKkEtAbXF7JEHELF4babgJxbtXRizQu31L/BXAW4lfw/Me
nonHztfxIfa0oZlbhdWRDmcoJb9NKNgCD9rPX2RRuxhmLFvO+Mn0LKnuYX3D3T/p
LoCSh4yDyH+YvWkpnxg+uvthlqeVaftWhqxCMxiqiyRA/hSrsc0KV/WwQzCh2tdm
BZMr3RZcAySP5WE96VoerQhbmNzxpUxcifh0MVRQnrQs4vN1cK4/gfgkDVscQvDp
ouBkZqhHH0Ps5qND/mx+d9DQSJP41+nZN/g3Snbb+5JBnAlnKmPvmP1SCA+YDu4G
65bPqgcEHCmt3ZJkMkcz/TCbBcyzbyL9NHALF4BGxVy6LT+nHGoxckdu5F8NT/9a
e5rr2n2ltrHN1cfqb9fx+2/2PVFFP15Y5en5S0uYXSSd7e92VrCJzWANh3e3Ltsv
gMxpTGlFn3lLR7A3um/Vrn6/mkmVfPmaFyv5UZhH2i7wVBPvrw4/uokRBdDIMDPD
COYHVJSHaw9LRAzVs4+c9peKZqoC5hrcEvL5H+kVIo8sB5b/mEfyCfchEqdsk9ZZ
z1ijpAU6DPnExOgSBHSD8C7Wt5EArj4eJu88mGj/qFqh8yxoFMhpsSeJ9Pgf4vn2
5/lDzyn7F6CKsh2+yvBiiMKwBA4s5+WnGoC+Uoxoav3dmTiBCisQnxdToN2FKKCS
Qs8j3Z1nHovZ7J3NK/fPIOa45uLq8YwUvn5P/s+Y/kfPGtU+3XTnDFIBHGmNNCsP
I5oS5pcszxogGopq6/iKLuOjkPE8qnw5yeYSNMyLmDOKPKfvX0RrZBwPPV8LmLNd
imsmSbkDUCXQEMqGAPuAqCJEYgyWEj+tNAw9TJixrzCVip7huh5wYD5QvR4Jqp6U
twtbLasl2xrwshc1X76hIvUpNzylqIfwqVDBThv3sZqr03JqsJKKq7gVhVJI60lS
HqSjA0gBYRm7pT5rsA3QtfzgN04j2Rfnlv++eOE/aai4J66LjqfSMA5dQTRqcPOC
OC8ymq3ELg7qnz/H9Iujalrx+cCA0laP5z7vThPdkUuyhd+BJg7PljVLG9agnZo8
2DRWeCc/nJ1LmK4v9gWwnWqZ4IUsutTBIWwxL2HbfhcME6rqL/U1MJgPXDr1ZMC7
EkpWKo0gVkDVqGqTt9AYXLPw2cpiHpJ+Tuitzl3RQz+KNq1DivjpFzel+hysidgX
SRW0fjHGcZAqXL/cwLTJmTMvFx1maENlxTysjwup7yxyAK7deIyZhfNQaKvGtKtB
PKfAt5HnYqIX6rgvVukLWgBNdGFZEm+OGTfab5941gYBM2f2RbPdb+5NNKeuQSHl
pjWbhKg6m9rhY4dWR0Y8U0MfDTnpOdA50I23AZEa5L2DAN+Iyk57CaP9Z5OrtEkg
F0l1mABXFZGqT00aD7r/yHtSX0DaG393G0RBtTsqMd57ZI7QxllmBODcG1S8C7g/
K4AthoB1QFAHmU2vJAODHnccHyxEpD7SY8CIqTEnuJXAmRfm2eELiHjneZkYAh3s
omldJRdV1zXF/dD6ysGRwZnPmtk995MaH8ULbVyUoAlC5buPA9/Tly8lWAcwmHdw
yc7CBgiXpOXCzOwXLgFs5QPynzu4Wx3L5odzgk9FdYIEowTmOQgeuaId6I8SY7gs
yWg8VMadmjotSxkLL2kuJuI/alMhxRuWmWc6yWts0Bo8uKWsgD3Xl/1UZxm7gxKv
tpL1QoB2rgJ9kSToR2pYVPZqGef1z5TxQ2SHNUWSMI6wRVoPUmp3kODqxAyDHB+e
ejGuqjwepLqYzsx2z0IvIIe/o9ehkFc+7YN8oqCRKqVuO4m6bZqaugIZtHfFe40b
dtQ27CeWYMMpk1YyuRHGjGMZVoyP5MxMp4UsUB4RTSULhyn18V2g0wgkjYwNWD3I
B4LlLb+FjgWMlSEPF5Q9FfcxD9bC7qE4ifuN9BOq6feD2zEKuSpaYGYqMiRwl66F
tf4W1GpEwtXtKXYoFZSLRh0lzvEK1A9mK93eLNbXT+US6SV5pPHUyPV8xHSVRTDC
5p9561rwaPzZR4pE9Y/RuMPugP890aqTvSd4uT4vLfZ//snLoLK0DjZRuGZXQ3zt
/cE21ErLgPL3QioG729OAQS1IV12l4p6psZH108rX7srj3hOEFe+NkD9lkgGI6G6
si1zm0dw55Sch/2VX8evUHJzhCQ0/3sFH8fKySCGVRShip6UgNoxG9Drs6e8GTFK
JhHDa02gIH5NTpERQOanRbMgJKBFJB6OfJnwRVyra6I=
`pragma protect end_protected
